��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����9�?5F{��`�!Fkh9�b@\1d��*��D�����=ˀݟ��"��i5�W	��*�)~��#����S�W�ܚԘ�d�hA�}1w1a]�b�x��zYP�C��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�m�F��������2�p��X^h��@��[iKd���3sΆ�@���e)r�atVƿ��ߨ��d�_5����J�&z�<�ܮU�eM�%��fG���z��k��X�D�]
�*�M�������q0JE�JߒH^7�8��=��l���@�@�^�+5�;�=�����M�1)�o.�5Y��9wgW>RŹv���bp�\�A"
���z'E�T_���9���*��O�N`T�(Z���y�dw1>ׇ�����x/���z��J�s" �*~
6�g���h��g�xH�>�^_T8��0��o����lz�b87�_�9��(�= ��_E�t&6EUX��cB䏱t��ԓ%y;gy�%����FH� �HwQ����y8�9�ʩ�瞺Wk�&V؎�#τ���q=�!?�Dc�ИI7��d5���i	�2��¼�s��퉶N �.t� �n<V
�*�niǛ"�ڀЄ��y�T� ׎�U��mb����?��T���$��ňE���,t4$A�@V׵�wY��`rP5�b��x�D����!��ɱ���y�k������gJ<��Ѥ�XA�jJ��R��s5"�����j��.�U�b��:�{Bhv�m0!���;�.��6LFe�;Z�v-;{�W���6}^$K�
��E=L�5��P�WgL��5͌<�+C�b�\�%�G��#K%���E(�*/c�A�_0y�_���x_L��*��8�����P��cJ;y��4��&��ykh)����\��f�;�ָJmp���J��CY#�Ȣ�M� G����#�{#��yzFU$��G4�%�����z�x�A*�6��m��+�z	�A�n)�����烉����Y�t�<d>Y�L6�L�!ZF�t�c��̍ Ԙ���"R�Xw\��++���,-��
��{��`~���Ub;��?���.`��Yl�_�4����F��Uvͦ� ��u�m\�/�B�U�Hs1�7/�J��gFg5s���Fp��Ӥ32�Wr���o]����[!�{�my7>?>[E�3��p/1�=���E����ڋ �����g�ʐ�2�"�sds��^lO&^Ќ��^�`z®z�%�O����Ȩk��ц�Gw�R�Y1I8U^��xG�����s=z���u�.,_0ܖ�L&s\~)�<�gDf� �\����eBѯ(=�7��������=�h�HN�>���Ȝ`៏#\��h�!������v�ʣ�����	�:�R}��0�@���-]Upeq���7���s�y����TWn���+�<�c��Y�}n��U�9F(�/ص`%̞-�l�Kvf��i��� 4��-{�EB-�4�μ�>cJ��[L�0��=��2���Ú���L8�����{�X'��(�*�`���i][,�NP�ş(%��\_����(�������
��,���նv�JΥ'�+�k0ʧQ�U��-N�n��WQ��x�@A�Z	
���d��T�룍�p6b���e �YGq16Zagt:�`�D
n�+QhZ���π�#�!�dUCz%�ɅG'_�$(��
[�<d%��n��N۷f���>�����*F�c�o|�"?@5b�X�J;s�g^�땅#A��֋��k`�H���tm(=u-���(r	�����3�ƃ� �Lv�o|��1��(���$��'�y!��ڧ���� %C��L�A�1I��,�� of����j�� �����esG^�.�*�0�0$�@zs�m,��$�K}"#��+4%�*%!åӻ�1�{�j��=o"�X���}HV]	z�U+�ˏ�Ϩ�v�A5_y�D�ƶE��p��S�Mx'&�q�:��X� ��-�Tg�<7�3K���"�!my��i`p�G�Th� �J����	�%�qH��`�dO��i�Q\�2���������U,g�-�C$M%�ҹa2Ƈ�����T�g�F#����]���'e�{a3��6���O������.U��e��I=1J ��W!u$Ӊ|�@�X��%xu=M,����0hv�Z���A�TH�dVVİ��\�jc]��Y�������rW��?�=���������䴃����e
��XwA` /#ˊ��Es�?�D���3�("�o;�r�t��'�2�A�),@��b'5���w8��gR*m��7�gCP�
�8������C�)zF��;%f���O[5�*��}x�sQ��:�g���!eN���4#�f�`�}��31O�`I%=�� �Ӱ�zc\la���H��>�㖨5��˹��/�B�g_�2 "�iMKtI�pTU@�
��$��j�'��j��;6����`� �U�=�C��^���������)�Tp!\xhY�~�y�Pdj�?Ձ��ɒ��{��.��*���!��j�F����D(��:A�P�1z�N�.=ݸ���@��*�v��S�P=�J���u���]cWe�ەLy�����Y��Z�I� �/����XA�H�{���������do �@w�[P����(Љn����G�����ʦ�9Y��������q�p�z0��z�f@��+3�2�G���Rϕ��a�\o�2jo��`��6W�l/�CK��X��?��O�굋�Hփ֬4���y��̈́� �y�o�K��>��F�M�������z~z�}��d�J��w��r;��h��]�Ve�a:i�.�J��2:�M���4�hU�BCnb��=�9}�>�N�R�&EN��	!��ъ~�SRgG�q_�z�+���C��w��a0�8 G}�q�!o�����ߖ�6y��� 6�,����X �e%��,{^���K���Բ�i�ӊ%?G[M ��������ɀ���~,3u7MS�Q ��+�Z,��e8�(k-Y�)���U7+��Jh���+��Ty���$��T9?���1w�
���d��������/���_F��l���W.u��K�hR�rG�Ž����wv�ۏ��؋��I�ЮrU�3w�H5��� ����Z�ώܳ�> a�3��6��0a�%D\萚���
��~���^9������%'a`�	>:ʏ�p���8Iܹf�yt#\��g��P�ã��b����f��H.�����g�Z��-��B�\�`��q�6fb���:�|���6���������'���	��I
jxI��^c�۝S��e��K�g4�Ŵ&�{DZ���\���Q��/f�>�|ߋuꩨ�,>�,Ք��=LR"��O��T#:��I=�Z��lM�E<D�Go<PRE%����L(LC��[��X%0:i3o�!�@It�(K��b��������S<P0R��7�큘�ma�f������;U�ۋ�:oOZ�,_-�����y8����8�ꛖ��'9:{g�0����	��&�)&��鵌�s#L/?�#ֶg �����zm����,r�	G�@iaA��1��#����r)k�h���p՜�,��т�tF7����w-�އh7�a���S��a�M�ʕ4���3��d$Q������zk���Ң~���ևr߭�vɴ)a�ˈ*6��&��g�G:_��	Z�:04���w��"�?���N�>:��O����,馺|׭�����a���>ᩓ���-Cv�#�n�A,F?��U�F��ؒVO�)�P�딃}5%J�
v �+q��)���s��et�@��4d��F�#d.�\^��{>�͎"D`�ټ��|�@�
E�D��#*|�(ԡ˶R�"�5���3�Dx�\i�g�Yg���`$Q�ުOv��ӏ���U�nE�y�FE'��Q�8/
����ys��n�CʩM�,��Xy�B��O1rJ�h��έ>W8[��ďm�+��g�����>�x�QV�HKJ��Iɜ�����7�7�5�� C�]C����ZUr�"`ؗ6��A��:"\���=�"D'��D�=�h���
4�H���T�/�@U){����}����nX=��m��8�ĩ��W������e+ɝI�3* ���H�W�iG|������@j@�Z����b��)�N��'��P�vX5�&a�����s8����6���k�%"0���¤L�2�2��������*V���7j�(�^���w�v�Va"#G��}�I�;\�����jb��#嘈Fx���\��{���ZheԔm�7�YVL��ǿ��l�
�6�X��X $?�xP6��W��g���dba���O:=3���%ų3Y��KDh׺��1��c#���zI�9Q��F�A���5�������-̶g!�X%Q0s	M?М�AO��M�+���t���
&z�`+ݽ�ٜ���.�@.��%!�7��2߮�!�s��=�SMک��0H��}����⩸z��݆��`��&�U�M�UJ�)^x�ۨ`�c�V�-�o8̭��WshX�@\���!��s�,����o�[u3���6�b��Pw��@5��� �oi��g,o��9*��x1z]Xﾃ�Uk'�����Y��k��D�!���;2����k���x��}G"��ѝRh����μ@�uu����!slF]� �/�H�� �cf�wje/rI֓�fW�����/}S�o'u��-�r�����d]V�e�j���mG��p�=��{񝘬^�ѹ���ƭu�W�K�UJx�
A�G?�?SQ㍳GJYߖY�l
y����|�)�;) �:�bk����( ORq���l,��a1�����v�D ��/5N,$�li�q��MZ�쏪�oT��L#�� QL��=!G27q��-}��Jf�D�H��^�g�GA���\�D����l63��P
p�Hy�5����$h��M�+ :*Hbj�� 5�3jGФ~�|&
mC� ����X����f��Ţ���w	#f}�5�y�Z��|��h�K��ݾѣ%7% �?�	�dS]�I׬H1L�QH�.�	�;��h��@��M��g.hT�`����j��H����kY��$�:���A���ƟUb]0��R,Q����QĦ����4B#�������I�|A�����@��j5
-BN�L�M{�fdS}-�DJ*A~A���
�k�{�Ҍ4o��}{�l�NT�
�X�䳕��S�Pg�r� �[!�fr�O�NQ{d6�r�g��U�ԋ��>CA��I�X��V�c�z<"^$r��������w�t�)�ݝ>�z'O�yX�uzF�"7�D��d0X�S�+���3�N�O�hI����U[�����l�����_�i���f���KcO��`�:(�l�[�#j�^y�ČW9��LJ�ռ�����	j�t�22��-�ڎ���IJy+^[����E����é��S����+�����ا�S���R�ͩf�(k���!z�j�T�~��}�F�hYHZq�<{��.�r�HjLz�
C���>�ofcəQ9A{���a�c;�O,x>��e4y��*p�{

�&x(}�T�6�.aQfΈ��z�`CN׵�w����a�,]&_��*�۔�� Ɣ��u�����MX�D���PWw�!��B�c3n-��I�lA��5��6�2�x��j�ꖍa���ɥ���#&$�'s�PDV5� �aw���Q��;3g�!' �
���L$�?I����R��P#��U�l�\B�+�]�����Q���Px���ț0�L���g��Ƽ�=�:�op����}�1�U��/X	�V�;��U�rE��ڴ�$Ʃ*=+�x�GϷ4����4��q�Ͱ>���)��t�!��3��>i[`9��*!S
2x^�p�Ǽ#�R�*�g�S���=�Jt��l4��}3��J�ͷ�	d������T�����b���l��Ǵ��ۊa#��7 Dy�:070�]ѵ��h�4S�'�J5A��&�S$Y9���8c$2�&X�}' Ҡ�؟���§�%�T̓~kZ�ؤ�3էݭ��do�7�;���6#>:��F��5������r�8Nā:9�}Ȍ�\�0|քC��8��'y��Y�e�ٱ��'ҧ0�;�!�ۢ�����5�y���6���ۛxw���q��9�(y�s�"\�y"��wt���:��2.���h�$ey$vNR[5d���b~H��(�����.�>i�ѱ��kq����M�`������)�9T���|WL)����YPQ�B3N
���r�}��{��/p����F�%e|ƍ�|1��JJ��N(�(]�#W>S"�a�=I8�J��������͔@�F���|Z��,p3�,@iT�LP�Y�-�3AE�xUr��e}��U�c��Ҵ�~�=>ٔ�f����m��	�y,zCC�*�M�/y<����nWό�&�)d�C%T��ў�?�	'`�+~���Ɔ��Ȅx5Ŵ*�=4��5�T�� �z!Ѭ�>�[oy�^�ƈ����=8v�g��s����I�5n#�
u׷�տ���9��0��Z��pF_����'�t�>��	G����c1{晕t�U�����>�4|�/��S�n��-��~PBő _h�&{�H������^&����r�M�������L� E�X<$~P�Ҙ�b|+S��N� [;�2�C\tڴȀf��n���.M$suzH5��<�D��D�~g��m�CC�s�=���L�h���L�N�3�o�w��x
�z&8�*Y�P�4񶛳c?�vUZ2sK�j��h�6�9�V���k�$�8�2د�N��gFu�HO�lH��T^9�Ӹ�џ�H�=��Ǧ�U\'��w[$�?���y��F����y�?N�H�����H	{�l9�[�����F��J0B�$`ڬ5C9�]5M�*�Bz�^�+�dD��}/��[�l��D/� ��|��H�m_�-�t��m':��L1DM��=da�y?L�'0 �^�y���w�����f��f}v;B��Z�E�S�CQ3�|��t���M4SA�A(ޖ�V�_��~~�f�5)>oU�&U������Rk�c��qI�:�t��Q����_5�N��|~?��<���E�"'{��{�2ԗI��Ju��d}���t�2D��Տ�V 1��1%�~PG\,J�Ol����a�;}�H�݇v�����R�œ�	�OͬAX�<CWo�>=�B�
�ns����#Y��i�.'-��%ǫ��_ S>b6φ�٠��O�lacG�����K����J����a̔c���2=�B�u�=�ޢ
	� �W��[�{z}��%����x��=�S^�c�i5����/Q)$�d��;����rBDi��������ܒ^�'�p6�V�f]2��[�0�T�)wV!m����-�?�=_�X������5H�Я{�._�2ӌ���h��N��Z�N7 �I����0��Q{18�PL��S7d�˰��[�M
��J[�qG�XN z�@�BU,3�뵇���0�:��܁˫���Z�u��	x�9{jwm{W�'���I]_b��$04a��I+K�Rm|Ӡ�0�fx<���˻��H���.��uH.�5���� �MA�|�R�`�i�;��c���M[�g�5����uqB�T���x��y4����R�?W!țU���������ۇFR�����:�S�0U���h���iM�:�vqc��(�Ϫ\�єM�!��^[��r�.�Ĕ�a�B
��0������+\.��� ��&�'����#к�K�D@c�8�~�[�y�fp�6c{l�\we�-�ڂ<�ɳL�^�2��_��N�.Д؃���?���2nR�}������=�c6q�R���$�p���^��T�a��hB�]w
Nj�o������-�?�Ǆu�f�fKsk�A�`��$�9-����-6�JK�6��~ �����̉��zFF�%���h`޻3��}(o:���:D4S?�hL
�q�A����o��`vw���b �ϫ'*%���^��>t�-���\���&֖̹Ŗ���f;m~iB��9C�H�����5�C�|`&°�ͱ<���XT�;�|��o��H=�嵒����E��?�f�%[zop��������i��`�T��[�Q�\hN�]U�NKq�����)�74|�$��j�gɌ��nZ������x������%�4Jq��̅����Y��97z%��'V=�Sox�3s�3CB���iô �2A��ړ����AN��9Md�H�T�Y{g1��?�w�_���.)sp�������W�hTөE��yD��w�]����~$Ιy��pz �H%�~mh�58�Brm"Ȳ@z��6����9��l4)ٽ�b3>��n�	}�#�.��tNz.ӿ�-z;�ڬ^��C�+����EZ(Ȯ�q�D���ȥ|����:�[3�������u�G�(�F��,9k>��Ђ�f����ek�>��}4�&��_Bbk΍�;2.���|�U�&�N��t�x=W�	5���z���Yi2Ḧ*O��>8�?���5RJ�&b(�ps��0��&#Xv�=eCK����)�W�,�ߴ��Z�ʃ�/)z��;�)�xˑx�4c�EU�s�#g�E�(��u�'%}f�ʕ�k�&�a9h�פ*}� �=���뤼:!KJ�g�I��+���ң<0���?B�Z��R>�w��Yv�u���������Ue� ������!%T	p�h���}�!����f����Ҭ���#�aV�XW�Y�^M����N���揾LV��ڸE6@�
r$:'�o��2�kO������eL8f���$e�} ��ƶ�X��q~Q�ғ3�X1�i0�R�{��a&���C*�ߘ��f��ބ��bj����	���CSx0��%�u��Y9U��i�F#5Ӎ6�K�d?��5�`޺۴c�U�%Le:.���?$�5�
�`�!���P��L�·�&gI`�2օf�<.���Ì�zQ�ƒ�J��c�АG94t���lX-ŉ?�*M��9N{��d[LA�%���퐲1��'�)�kp5dYU ���K�'����<���re�c-|��1h��:�F��C]2XA�2Ž=��Oz������<�5Q�h�C��L�VR��'*cQ.[c�$2.�\����cb�`����I�=������7�&���}y<R��~}�C�V�ڬJ����X+Ar��!
%�]a���|�(�sJ�%?z%�nA�2�_��G.��
�SQ#�Y�V�*p�ݣ
{���F\H(��6;���^��l�0��;G/�S�;�*�����=]���O�G�޼T���A���~�n�<����Ou���נ�+�3
/+��,t8�x�z�X��
����C�+�	�i�"�n}:��@ވ�܆I��
/�YC��9����g�w��E��~�h"f`��䯕䐊�-����\K�,J�mVO}�#����YjW���=
�2�:��-��Ő5(��^�y�~EhD��a��Qv�@��i�1��t+Ѡ^���i�s��D�y� ��xTkP*��F^l����ں$EWq�冏��S�eJr��M�GƲ"dӝ�6/a(}�F;�W��s.Fk_���`	���..���V�%��O��3W�orF���Q1-)V�.j��/D3"?i�>��U�pK�7B��*��H$t��	�)�����8�y��E�0���$v>�&��q��L��&ὗ�{�O�(�^��������Ǉ���7����.!�s=�/�/
\��U^��:E[tA�M
�C�^���7X���ڣ�"s��!+b_h�D������V1L 5k���Y��6~.�Ӈ���|�|�8�г�f��L��z>��N͜=M�3� ~�r1�ꏈ� �-���o��5EA,r8c�O��ۤ�&�5�]l�{t�զ��r���.L�>�(��p�cS�K�buh�N�����Fg�b� b���+�)O�)��>w��iF���MJ�C�J�?�N���p�<�����GX_��u�g��
k�"�z"�Z�����3�̣ �	_%��L�]�腚�*,n�rUR�|�\�EC-χr9Ǯ�� +>NZ�� 2���g��\�k�	�@
f1�q������c��<O�%'f�V�-����!��2����K�;���@S)�և��z��}�&v���6ZO�~I&����
s�#��^��wn�c��/��^�i��&�u����XS�72�'�Ł�d�o;��&����qN�[Jֻ����@3���BLS<�M��q��74B�o��v$��Y�3�Ah��,��0#�K��"�)@�Z�f�A�1�}�iT~��
y(��f��$q�a�OR�K-#ƾK��xy���s�9��,sc�J�`��-)Jn��7i�8<�����᪜���5[�g6b�aV�	&��O�cx�@<�7��}Ld�s|���N�e��P�.ݘ��1[�ϘZP
�is��!'�+t����Za6��\�����I������6���q�(f�sqCL�uTM�������_���=R���bf�Y����c�1�2H_��d���ޱ�ɓ��m���6���Lv~�Iߵ3��x��]?������)�w�����Q�r�H��g�Zz�];�e),S��$��Ki\��63Z(ҥ�-\O��Wg��B4Ez�)k��5���䴊ۥ%�St��@�E�}��H9�����!�>?o����?1�hċ�3�ڔ�l�u�� ����AL�H��^g�������/����#�|	��93D��7+��m[�C��wDC��X�jH_�r�~�3!euv����k�q9�0zaՅrҺ���-�@�g��J������V�r4�C�hU�tqH	B	5�����}��;۫�F������En�SE�S��ܛh��P��i����g��Զj�%B]E�A>	�\� ������Yco��w��9rems�,��ϹN,d�p�"���f��Ќ?��]�I�v/�2�`n��a�8bDy�w%��,v<��\|��G�d^��3�
����b"��s��ˢ�OW�9KR����˘����cL��h-B#�^��bQ{�mF��X������{����F��U�c��%g�Ц��}bʜ�zA�<Y�֌T��K��Dt�4�$�"G�������ӝ���mw����:��֋o�ݭ��X��G} N:z���_O#b�X�=�5����->)�)�` HE����'H}�u�/l��cC ,�`�	�b�S��D�!�u�b�6I�a��N&�!(�}����3��ԺX$澜#���x���O�.�k`�G P��*rG_s�=��w����6ՉY
Qף��m��Vа�M�6�);|.�h�ណN�x�2r(:�8�z,���pz���S�;n�
�� v2�y����n%�Ȇ�,��K/�����lJ�"�"l��1tr�p�<^�U��w���������{Z�N|�)���a��.�:)�˹M탌�i�����Hx�g��lW�7�6��"MD�hw��X��#�8�j�W�9k�Y��r-�R� W�Qa�11T7��}w6H��.�u7WC�Xm·��J���i�V�S �<�̉C���N�A���;g���>��?��
����c>���������%uWxx�xQ�"T6&�:�f�N`3Lh�6�T��c{y�S���_R-~id�!
��_�m�/�yf�[dז���%��
�0���<��q�	����br�j��:j�K������,�Z(�J	��Rt%��Y�HG���������ԣ��hYU��7���H�wbm�W;"��Eb���x�5��,&$������ڹ�Ě����.4W@�i�!HP��9F�a�{l'�:�@�J��	��5ɪ�>�;7��j�q8?"��K[�Ъj䝃���Uɞ��l�{ w����^�G�f qj�tj��]Λ��i 8{Hk��~k s�˄�i"3��U��]ΰaG�V���a�~)��?����=��:v<� ���i�k6.rQ+㊁2�����ZW���;o��4�^������&eƢ<�ق�m$���Y�c��5�A���u��w�}���?y��A@�t���#K镸�����O*�J���5�Y�/X���V{Y��V�t��1,��)Ǘ����&��C�Lz�j6:(�6Yֺh�f���M0�����@*xzp�Bi3��<y��a�f���5��0�^���}�Ю��c2��� ���Q�ǰ�v�����|�
�(��_I(��Z�J�O�kN��m�!��Ko�.x������a�E(�w���vZ��g(F�5�\�@�&C�3J��]�g��``$;7�3������G`$XQ󝙕��l�iqG��a
fo����Pi�����g$�VusL��<����!�	������f�額�f*��	Ϲ{��Qfx�2ij���y��#�F@�N���6�ӝ��#B8�נz��
����j�V�;NT�Փᘡ��THdH'�"D�^-��:��(��w.�v�pk��xʠ��>:*�����q�ۻEǅt��"lx��/u���,�ޟ�h`�T:8�!�5�3�U�'�<��p�� {>�Jl��g���]�g$�v�@��y���#�jw#�ж�<�{�e e��O�]&���$0�i��oRk��մ
)�cVԄ���WU_5V�NW+��l�>�{Qꛃ�yC���7;��ۋY~xq3*-
�]�bn����+z���-�2n����&/���2��6��rE �R�d�7k(ZO�wx֖@Χ�l�����v����G٧蔫ь�UҼiɷwGo�K��6�9cA��-|��ag2�f@�����k2qk4�Dc~���K�`�.�F?G%tM".�MGԡ�"����:�� z���Y;�'���^�h�Sz���?����4�w��{�}�CN��TI{���ޡe�e'[%�jTCW���-��ǂ���20�����̲��m���w0�Fܘ5��gq/��^�n�8:K���o�2ϯ��s��S9%�����A)��ԝb^�c�ҊK��Ц��o]��nr�5���콺����s��[�LM%��3,�����v���ۊ>H��!��^0�Ҹ�x�>�r��_Wi&��1��|[�R\F�Ra(���屪kWd+����l{�떇af:ڗ+lo��_fh�W�0��F���Bbe)�[aY�Y�,"P�#�Wx�lu𱼎MJ� �C���|�g��ס���`�cz�3�*5���=���Ve��Y$�B��u�΢P-M��m�3Z�b`�J2�T�j�,1������(��L�GP���a����3�	���'Kl0?u9 �E�ۏg�}��v�R���u���HGZ.��1��y��sw2�@6�߅�poq�*���Q���lY��֟
��ar�<��&���n�quNZ���]y�I+P�_�Dy���O^G,F��S�/��%R7�/9��F�z��nnU�??(V��l8�e���4]���JLF*9���]�YQ���-$���DE���2�ٛYz�����YJ��4�G�f�!�534�#=�3�\ᅳp�*=�?}�Lz���5��j��#�!�.L*��/���8殿�Q�<�ϝ���0���r��1��������5R$ Ԡ�����V�JA���-���������9��mЏ(��!o�>�e��"�ɖ��v����̾�0���?�@�p� ��^7�D���2���F=��/!D1AV�|)�;��ddރw� -�dw��u0ߕ�"Sd�Rm �$c�t�£G�ŋ��hk��a��Jtb��a�l_��@�r��r��)^c�B4b� :Ɗ{~\�/D�t�r�I �%**w�V����3��y��p�.�j���S�7���Y3 ^�r1#tfM[P/�{�F�D0�-�MF��$��1��B���	)�mQc*���(Z@���&q� �(�V���)_�+e``��]�>��ۓ,ꃆPW�j�+���:�f, �h��5�b�TW<v�(�kl�
ڶ�h;I͟��i��	�C}ߋ���=�p�d���о������r����wh�pߢ?�%��4���-�*ނ�-� &����#�,H����;�>~�6-�K8ό�]R[d*�x��c%u��f���c~��|�i3�qF�U4���Ν�'���.ef�$�rq�l��h��؝%��fё���N�J搼��\�z���
c���+�TJ������x�[2BJǮ���W�E2Rb�J¶�1I��PR�3}�4�����,V��/���7o�]&!�yW��+�����m[c����Ӑ�`����.���I�q�[吀���<���*��Y�k�K}��n��a,6�Y��9I�&�"kD}T-g�in�!��:�㕺���v�D7���^���Y6f���fP�Ķ�����i��V,����椂�I;�>Y)����D#�ٞ����>�������n����?���E�����u��$4����c���gtM ����{w2�=Ȗ�g��0�t�p�*������O5Ue�@d�/oC���G�#
=���Cҗn:8�%g��	ǁ겼�Y�Qm��%��O��埫���IK�hJMK���?���]�����J+�6(��!�Wmy��{�!��Ɍ���	1XT�ۄ�<Ո/Rb�A>�E��}��0�P�`�?�d��y�0���,.o}������y����'���_�z��� P��ɻ!�Yj�,���uz��F*k�P�p}�9]��9��P~���m���'�ĝWlx���32�Qt63C��$�>�h��[�ˍw�Ht�=�|祺���|����d��Y����[����n�;)@J��p�ٱP�I<��X-p��MI�6�F��^�CȈw������	'��VP�3�G��p?G<��CQ��n��b�a��A]5��X�ﯨ�w��.N��1�fZ�S�bi��׌�p�8�eˍ55��[U�	�H�|̾Z>У�o��6F7��:������N��t�ȵ�H� ;cY�nȨ�a��Wq~�F��i�1��@����m�p�3k��T���P0M���<�?���O.�9ʉc�B��}�>&� �#��5EGOT�Y���=�}	;!�J�g��Gi2��Ǿo1�_�l�2_���By�F4��#��l��l�?��=8�K8��7�5��*N!6��ǡf���.o+��a�Υaň8Q�ieh{;P�n�@�%�g�Z�H�"��U����j_�y�^g\f��j�oh�N��s!h��w9��Y�o���b;|�_MUt�����)���j�j�H���J��^�1�m/�*!�4P�U䎷�S높J�n.��=�P�zI�J��sIގm�)/���~g�`��C���|�c����I�0%�6�J1��)x���'K�۸§Z�:S��U���M�~�=ɧ�Ŀч�p�P�/�mu�
KJ1�T�$�$�����?��J8�E�α*�	��L*f�Ҭ�)�(�H~ ����Eօ�2wy�,^+��=�����]�)F�m���[�{�wÉ�_�Ns�qW}b�����F��wX��W
�A#�?�ᛡqT�n ��e�\��
*Ă��?P�}�D�'	�գ�8��Ye���$��X�E�M����$�[Z=��0���<��?���l蘍��H�9#�<�� ��0�����|>����o�'�<��<�����cc�e�h�|�$����2�lTF��x93�t�'�.;�����x�ϊ}�I� c�VϜ��k4���`6�&�^Y�T}k����[Ŧp2�-����䈷1�1o�Z@�u�Z���-�.y<
>�-L������̦�fo��aA▏�h��Z2��p$�yC^Xʃ[3"AhD��,����p:���Vz�`ըYS�R.���U�ڃ|
��Hb۳�����hx�,{��<K������(��+B���3�r�=Q�s�K,�o��w�;PoCɷU�Q	Ӂ�_��e[���id�.�+����Jڇ{P��i���>N�m�=MH͟�Wud|��z���YUZ-9��nrbyc�2��z���Գ)�[�#��Zz~���'J�U�pt����~��KjUTL�Њ���o�[�尶��Q�K=2Q�U����n�dT���金qd�:�`ވ��>� ͂1�5^��D�ͣF38� a�]�(J�0��
44��pQ@"jr�R����,�C�Jk�*b��HȮ���f$��d	�`9��XYo�9��Y�t�� 4:7
^=j�taLWG09�S=��S������0�8X�6o��u�����#y�>T�	���a��l�c�{`5��;������YZW
��r��TX�������8$��~�L|�	>���K`ϕ��1�\�2�kۍ5 ��PT�ơ��٭�	-�?��[�P��mC���k�V��J����W �|܈!�;>�l�v_�6s~[(~q'������J�ƺn �7��z���j<A����yh�M�J�4�����U��S�:�uW��,�[��'�EG,�w��k`�;�[��'��6��.J��A�G9��8��l�})r��R��fj�v_'��V�NV����\�'O-��}S<�d����0?r8�ܙ�,�O=8�qY�5�; �*�?�j+�Pl�ܕ�w�Ҹ�
��]�=[Ou����W�g�~��z�`w�"�gᆉ-��i�&{�zU�\_�LeeR%=&�����z��An��2d3���=)ӷ���c&��S�[�γ�޸�(��"3���m�2!Z�O�FVG��f�1��+�V14C�<�����f���Zpge�ME��8Q^$I��������?+I�1�������E�$��:�Qh�4�%	��8F�7
@�T]�Y!��\�C�HR)�ݳ�.�p���s�Uw,U1Li��jv9�<���1E��'4�֗�Ļ�O��ˡ+��80!�N�k\x�8G��o��W�<|�1���E�$-�K�}e�ѷ����3{�MS��G�3-��
V�����ۢi��X.�<�xkѿPrl"�{f���=�5]�A�q�"�ӳ�>�馭�A�!���"߹��@nl �|�'�a���*�y3d�A��F��L�S�t��Ż�vg��->�PO�z�8-�����WX�x��
�b��� �W�lb�%��n�/�k��e�����C�t
+���#hcy=Z�c��eȶ���I?3�{�&�������M;��6φ0�����_�c۸K&5%R'��q��6��\��fE���L�3s��cx�)�_�����#�<���Y[~xaj�Y�W�%:U3���>)	���]�F�d.!�xڥ�D�\�c�lX�N�J;�G_p�e����xA�~�R�^��Z����bΓVg�_~í�y,n��F\�
���0^��s�]<�\ P�;���He����;sA2T�nnt�
�� 9>�.n�xB�j
��e#�j�q�#SL���7A
{}�L�[�׬��?ᨼ���
k����C�j�`mCd7E��C�����A2\!y����]frQ�(�j�nu������F��:Ӱ�Z/��M��N�]׌���mKl�_� �1bAs���ǥu������}��F���#��O
�8(�5�����k��'�Y� ݒS�G�>q�{�P"q��1�B�2H&[�;��Z&">S���*�������c�O?�}�c�4����N֏'j7����Ludj�4�!�pK�U�%T�b��~"P�yB� ��Cd���Y6�j���o`��חE>$�5�T�zn��LZ��o��S= �A)7��.2�6u[/�Q��i<�:��M�Y/Gx�xD�����Y%� 0�/חl�ޛG��ߺ�_uV�u�D�g��Ba���?�̆y<M��~�~�tC�>���R� ��\�ڻ�)�qE&�B0���O��n'sd' �m$v�m3)�lHD��˪b~��:ElUlsf2+KO@��g#�ߒ[�*�{fd�rH;��"����M *���wh�Q'�C��ۅ���z��%��Sj�TP�\b��,�ӏA	��_�˂o��c�ĉg<�|w$�����	 O�+t���5i3F�,��,��-��y9�L�� �knE*�9DDdgs�Y�z� ������#g��Ck�Q���7�[,SL��f3Ɉ����U`�l��])+�j/�}3!��9#i��K)nCU'�J����t"�f=�J��wO��<��Uh)���B��W��ػL�������H��h�U�bT5�z� �^�w����~CW������J��@���e*|lޣ�Ԣ� �a��#Xn;8��b�����^�UQ)V�k  �Ͷ	�(U�'i
E�c�`�3�'l��Q-/����b�S�X�g���j�4P����s^�/(r���{L����@�G�� [�>0P�'.o���5F��j�}��w�ʺ@��mdM�]rW��S�NM�m��*J�J-�s�d\���~�6�k��_n��\��F�f&�Hs;S2�N\Χ��$�,� �5������i��GM��Ȝ� {ZTM)�(/�����Lw`Qr��<)�	<Lj	���_�+��>
��1�Ƴ�e ��ᯜ��9�����0)I� �u��G����k�R��B>�7�����$��FA�m������y}f�iU�~�)ķ�koV~VZZ<�{��x���M�Bk���kNF�(BH����b��駂3�ۯt�Y/�M��&p?����a�TZ�`��E؂O���׽u�?�(e��I��^�jQ|#)J����)�(��w�;��Ю�0At� 낯���
�u1��4�����F�8�菐Q�s����]�My��mVJ��޶�U$�~ [�(��^��H�{"�=�ۖgO�W���ft*����$Wn�``H�Ϡ�6���͸����OfD��\?es��/*+YN�)<�>��ſ����� Z�^�τB���TY'�o�A�-�#�*T�8s�Z��ȍ�=J}�	B�~4��]�%tڼ'����hW��qX��B��/�� ���C�h�QB!�a9j�)����c�U8�a򋊟[Is%�BNړ�r���}�nF�t�Upۯ�p�f�\r�*:'YB�V$����)@��@�]ϻl1��aDvOՕ^	�H/^"��Q���N@Őb�-��,���Ɍ:`�k��X:=K�u?�UG��#�=2ҟ�4[��=��Jq��
��ǉ�>�X�o����N;?Ւ��^�|����om6x���-fc��K�AYIj��^@j�7u�g�f<EƱuF=�����w��A�^��kh�~UK&.�@���E�$G���"��s9<�|@	^�Fp�>2� ���0����U���|ԄP=�g$���@+w'���pOM�	�OǢ�D�1f�����'~�eY��4YE��e*�$٭@b��2����:�8�Z'�p���&s�7'E p�*J"z�}��D-�D@s�'H�kiQ�a��.��3�� y�ʇ�$>��'ӊLv�խ�ǭ��L��t3Ӵ�W_�����J�O�ԥ�O;��f�qЏ<��>�DU��Vx\uq��Z�����|+8��ˬ�6]�,E[^�C�hK��\����^�짤8(��hi��<&�UnhB�d�ox�N���sq�3)�Bؐq��U���l)RG�ܮ���?��g�j�.(���#���l'r��_1r��Yv,X�PU���)S%�-�쏥ܦ)F��
ϼ
�p變ß�@O�LaM5H'a���`��-z��BL
�/�SS#�9�b��e�%�L�{���u�
4�S��p� aJ�� JE��ip�������Ud�{SP�5�vɪ�$~��PY�I\P
�����F���k�H8��lh�z�Ƣ�^�1ǫp Nr���~AC�9;����S#򘼍>��K�f4.v\�Y����*�?MD>����_R�{�Y�#�{l�	|@�Yܰlp�<B�V��[ݚN,�^�8%&��~c&�;3��(�����We�|���g�ܓ�ہ��9���澇��l7[X�M	�]&�V{a�~�@�b�I��L� ��7/}�,��p�=�@Va�^�	3���g޲Q���8o���@�'*#�-k.0	���de��ԹZ�<{"lA��!��� �Ap��P�8���zN�F�N!������QÁM<��w�%��
��ۮ�n���w.���vI�;B̹H�S��&qɮ<Tˁi�Ny�g�>���b|Z&4d��Ӱ�x��8�[%7�~����Sۜ)l��<� ��HG�]��<����Dsl��ݏ�`7<՗@�8�HZ'S�4hX*X��f�� �P�~8 �4I��0U���Ȉ�V�t	E���v`�&w�L�%�/����)�
�!��<M�+�����:�nKE7��.���`�;"�@u<��jGoz:���pU	NT���\;�l��~'�,��<g����פ�WN�6��:����7Պ)z�83���.L�>��*�^�����b� �<��L�)z����oi�Bڮ�t�^�Ŭb��X^ޯi
�w]�e{./V����i`:Q~GM$⾧����t@�s���Ȭ"c��OW�% ��':�S�	�����݆hO���W⦈�L�4"u���ûQ�>��j�Oo���{��!����m5�Ҙ�/rz*�8�A꾖2������O�3K�g75���b�ҕ+�J�R ���^�p:�)�"(*��
�CY+��(��(t��r"�7.b���������ğa�=L~���;){��+0�˩C)��ﺟ~ŷ�DK�5S#���j�����(]�7Ӆq��߶1�G����b-/Q�ŵ�+�7MC�����>��GO��=�%��g�jJ\�D�� c�s�&j0�h���t	�mc���j�I E��g�D��_1y>�ؗ;~D�U���,���?�',6�
e���䵡�]�:S�EFϹ4��>Ø ��J��(�4,�� ���7xΤ|M90&22cq���M9�2m���K�L�8𬘍R~�1w���⺁�o}
'%�1�~�q����`PH�l�X�%�ϋ�$Iq
ˡ���I�nl��S.l�����f\��~"64a�Y�0����r��E��eH�^�A�<̋!��F�p�P&a2l��	O&��E�R� ��cТBko����S�j,5�0N3�}��j>�]�2���h�tsѮ[M�q�¾x�����gt���Qu�=� m�֒!zwRu��v�b�����`&	��=��n��	3�]��L���y:�����n���A�1�4Yɵ���V���ٓ�r�k����H	��0D�6�� �]�tJ4�M��O-���GH�Q�g�Dz2���&�yyJ�����Qc38&�4huy�gKj��3��=똛�@�A�x��"&0���w��+� Ά��%�w�f!k�V�~|H�j| CJ�R%�9��
�,��/#ɪ��3cz$$O�O^}B��$G���g,�����o'�ŠG�Q)�����.I������J{�bE�M�`��5Y?Տ�����=z�]H,�����k?ۀ��s�����V��L�}�vZG)���禝�:�� �ӺL�Z�v-&C.�7�v\M%Ha~a	�w2�#����D�zQRɲU=��$�$�O[j�b�ED�op�VC�m��l=��Yzχ����~y���7u�~g�E~�{�eA��7�t[G���u�Ir��O�ޔ����P-/��v��h�٩�X�?
�E��F��J<V>�&���E%,�/|�LGk�����Cƃ�����)��M��FQ����m��ݟ�-HԬ�X�����7AGY9��&�Cb�Z��s��un��IRB�����
(��{A�W�Y]w5z�{mk�lӠ�a��,̳�aY�/��k�=�6^K�=j�t�Z�t�)a���t>?���];��⳾�i|����R�RV�(zp�-_�o����5���a�&y�]� ۝]_r�a&i"Iw�h�(���(�7^�7:k����#�,z3�lFܭXxS�������o/X��y���R�MB��N�y���
ʃdߍ�.<b�C����/�-}[ �WIB��K�>�U�ѭwSR7�#�3� 6-���s���h��]���էQ%s��h�:��7{2�&��?�R�cr�ڇ@\���Z��������i�Vބڿt�ZZ9#E�O(�@��F���~����YOR� �"�ViA�s�A�U�|]4�P��$GR�sbo�5�������%m��EN׃&��Q������Z �?�?�%^-v����@�q)��R�i�3gg��&��tR�%�W��]+8�=����{�9���L�qԞ�@����&B���2����v�n=�v�w�J�M�Ŭ�����>��a�,��81/��bYs9h�rضE�tg�q��%��7�B�MG!��]"�-?yG���|�gG�Y��/�묄�Ĕ�)[c󟏓�I��NgT?�`��}��v��`���s��Z@�/{�u�9*����1{�����.,�o��F�~̀�{�u�J���Gӽ��6L?��ENO����և�0�e*r�E�l���n�%�+��b)�[%���#�l%A	 �DD�$w*P�b/zz�s����WZž64�t���-H��JPͭ�e;�̆cܧTM����C�sށ������������HڪkuE�:']1l�k��ۭ��_�A�%I8�;�ֹe^��f�[����������|�	ή
���L�$�8e�O�{���ݐM���>H^���ET"�Ɯ= Lq)?'m4'�K��sT�V�QyV[��߬�g��Უ���uz؉����/�b-��0������&K��jeS����5��=�^��
RN���Ss��~n���Cv-#��>	C�[��)��v���m��:x־;T�5ʅpio#��oy��㷧4߷Q!o�eB��p�|�Y�����܍N/ԫ1��W��.�U��Ocu��RX��ï]*JT4�O�a��+aU�����<잛E��n7>x�<v�0�	aR0����F7��7�wI|��+8;1@ql�G:޻���jW�ju�o�1<@26��-�е�����ƨ��*>4|?,�f�������	����.n �f�� ۣ�������4D��g>�<�V�/�$�`e�v�	����E�>δ���FǐD��`hVcr3��2�a�i��:���./	Ue�~
�0�O�/�K�h��s���?\����!���azME����G�+9�1Dc�a��/"0��>��;�l�3�9C�Qd�KV|�N_;@dY�T\�
8���A��$f�����!�}x$�x�^皛�cx�%�-�|F{�m���x�����i�h[`�i�p�G�ƫ�YY�����i�)�X�����*�1(F��sBF�}��ެ�_��ܦc��tb��H��h�x�zuL)��HދQ;�&ny��Jd9# ���D��ᇇӣ1&:$�	�{�x��T!2�����ِ2N��F|�!�!��Z��}%O1���I�<Y�7h�������ZK���Ѱp��)�xd6-'��$v��^������&��&;a���
�I��:������ڤ�b9'��4��؜tV����6|�oQ�fj(p��!o�z��S|��A�󤕮��f��������uă�h��s��_佼�z��jOw�Y1?Z9�b��% ����u;��#f?1��C�2BO�3�u�X:����k�8��6Ps>�!
l�� mf~!K��^/N�X� 0��M�@���
V_=���]�B��7n��`IwiЈ�,�(R�9f�'cJ�B�C-����5S̨L���������mD���D���}%�_Ը�yJ81d�O���%�p��
��>����f{P!wd�<0��y�b�!����)Ht.9�tDи����5�~c���%Bg��S����T�n�s;���]$R�~�w��WK16�>r4Y�݋`9��p
��cX/eU�?�\l&��1-!X%x&D�^�G5˘t0p]��8C@�+m~�-���[H;rĖ�.�n3������p	��nU��o�Z>e�Z^�o���ؖ��qz�[�3K��k�v��C��]s����
����ڑ�ֶ��vxM��4�'�_�C�6� ֬$M��t�`�/�?����h�S��gȘ��i~֐Y��*�$�ʃz��Q<�>e�*8J�4=C��ӊ�9/޶Cn�����x�����݈a�[c$�c���5�3��[� r9�1*#�E�� w���������=Y�T�ji�	��稙��t˱{?L�p��E�`�`�w�#4L�J�&�K�<����B����������`���m2a�b���Θ6���O�0wM�^���p5�7����.1t6G�`)-]��z8T߹�����`j"�0��K�D9�uk2�x���l�+x�{%�bScD�i˦�������$Pa�=Bh��{�iFum
�cl�[/4���Uc0��dH�Kk��nǔ�z�H�<�7wmrz_>�k��!�^�G(?���}��1'��]�^�cA���5	}B�����)�w��S���#6 ��g�ٌB��6�W���zZ��.��KS�>ơYyt�; l��Z�P��n��=�b)��-E�u��p]�m�U��h��!F(�j��\v~����*D��2��V�3�e�/0���?Z���Jz8/-,��&�dY�]�fţ��K�U��g����������c!f�)�hZ���8J��'��{>jY��	
�N�L���3bXG��W"�t��`f-��s�/����Ԣ��WK �yҼ�ǋU�e�8r�����%`E��?K���lf�)��6&�QBJ)�K�����pa�EH��.L��Z��5QJ��(W���k�6zw9�שf���}c��g�J���duiGS�[�5��)�›y�BfI�bb����X�|��n��n�+s+e����v���U)��c�r�5���m��҇�}O�,'e�9����yZ�B��춈�%x�`xUн
(ް��
��[��w+Ԣ����6:{���
D�]%wF��~A��([�ߒ�4@B�WF�����M40�G�ZN��jr��r_i�FE6|{�M~U�9� �,��g�, K�΅��S��DIy~�q�zs�8i�`�H9�lu�CG�QŘ��v�'	Ͷ����om )&��)u.1U�Y6hl��Dd�}��s��*��m��u�S	:�m��J�U�=ץ�LH�.)�`u�c-�&��kڸ��?���]�wN`
���:�1��'�oF��D�5����߻�DZ��Ƶ�!W����^o�"9�i��_��j�F$5��~�@�W��ǃ�?��ڕ�8�~��nk�c���}����:D�}swm��B>`V_]�y?��!ikC4B+��MD���C��{�u��L`;Ǆ_]��b�-������D����c���B�>���+:c�86�~Fs!$_x�6Ҳb�#��o:��R�;��f_��(z����ap$-b&�P�N���{�e�K|�j+�- ���1�E(3W�7�Oɧ+D�~ޜ	|\��Q"��f�
�@�^����,I
 �d\�`Ǯ����0�ߵ�0�������I	���u�E;�#mV���8|>`�Ai�q`"|�"2A#Ρ�X����ܵ��N*�`+�4寥\�I�4rBD9��WO���X�Џk � }E��6�H�vXr��
��j�mRI]ɒ���,\�,IZ���n��Fc�Y�fA�< fX�6j4�Gh���%Գie��mF�(~�L��/��Iܧ��sr�6��>����C�LX-��o9�h�G�[C�"���*G���oKO.Y�D���Щp�M(��3������JM%A�tϲDb�\	�q|�:��"������Q����V����:�p�U~�p��m؈.�e ���e��L���h��˓�®�7C������?b�2�:0AT��4�|�l`Z�:տ�P͌YAT��ߺd2=�9)�ۮյ���#{>�M��6�e�*0��5���Ct��a:G��])�H�)zmY
��w�bc, �@3��@`��s3�ط���]�>r�[2���s0�H�?��82���#�*,���&�[>/�>)|�6����_3��v�׉*
�F\za�[����;�����fb��������zp���K5nW���ػW�.BH���v5�Y�|����ǲ�S�����q���rw��u��ڔ`�ڛ���]�ן�
Q'�	"��[���p�WÏ��Jp�_������O�+Lh��*��K��IK�""��?��Y.�޴~������$��%#� ��ƕ��e:8K��7`�s7U7SV��K��A�:X��Hs^��C��ط�t�9 ��ڜo���6��Q(�y���u�C���'� ���k[�{r��i+X����-&�q�3��T�n�B?�1[�6���ym�wǩ��p�ݒB��ax��~�0�v��H)ˬ����QLk(��#�4s�� ��g�z��.B��l�aw^�C0��0X��� ����J�	�i��*q� B�C~ϗ3;��n=#c�u�����%W�0�f�9�x�C�i͏��}#e�M�2.�܃���������I��-���	|�Ø�]��]��υ*g���G3�fD�_gO���k��
P��O/�c����{\�|Cui���`��X6##�,]�
D2*[xI���F);v&) ����O[A�d�dJ��}4\������<���O���s������X~<`[D[1UG�Qc�(����+���bHʪg۞���<{i��nL0qy�~A-E��_���r^Ν$�H,J��3y��[Κ�Y�Á���%W�%p�SK�����ο�()�/���\��?�׮��y����x·�C��B��b��dQ[ �2*`�j�$��·��:��,�Mf7�*/M~B�;�6ݫ��̩�^H�|Q��Jx�����d|Lv8��}b��Np�{:׹�~�^o�r!���q�B�ǰ7O1�����CR��>���=��W��_k/���X�%�����+jጲ����s��X�T<�;��R%#},7����'W;w���L���}6��:A~dk%$;˨��w%�|P�����^|���(����f�v��
z��=i�JO ���vXg�M��Q���DjV�G ]ex&�٬�E=3ɡ������7��Xpz<�G�V����k�a8�y�>35��>�ZAz�^g�?���1�;�z����B��!�YW�ځFR�Z4X�g|o����iA�!�"�b�,Su�Q�h���dyTۄ%��A�i�Kfc�� ���8��܍v����]v`���Ǝ��W���z��.���Y";Q���������D%�di�̷)���x�]��ui< �D���p:R�3�BRM��x���%K�
�{9���,�+Ε��[+�#�Cg�b�ǎ'�
�^���P/�84�	x�D���I�u�ښ���Ķ��,��:Q�,ڦ,%��7�Kp��w�*MTc��)e�1�uH� �&vxL�Fs·�̎�Xi��<H~K�ʧ>������&���̱��[u����(b�_�U�ܗ���ف�����R��I���o����)�0I�����<k�*�l*+�2�b����'1�]�T��+�O�����������n��x���$�y��E���! �g�h�DD?��"]x���m�n�4�֗�ce-��	v�Ց�K����"�do����C!V1��~e�~c��� ��� �%j��
l|�ь�}� �^����R%���g������(��n�J��4t���Q`���&���U��j�ڸ�0��J���[�*�y�e��们���A >O�ߐ�Ƭv�$���]�%v#x����ͳ ó8ģ��t��m560E+;���!�-{8U��l(�&��I�(�W��������>y��}���H����s����oݕi��Bx�#H$�D��Վ*Ӹ]�U+��߽3"��a�&�|H�e�\���H�ۏ-��	��qC��'%5x|�5 �C�~O��{T��70�e�O-Y��Ww̽vdC3����3Y�����������0>��B��9�%ts6/�U	���mʃ3�c"�'��>�m�W���//�* �#�.�U��2���A��R�C� ��ͦ0�+j@���yYN'��I&z�{,8z#�ګc�}�k�O C���a0j𐦰��]��V
5�(�9H�`\vR��Oo\DhX�]�R���dš�MW�0;�"H$�+�A�ΜI��ΐU�j�B��2nސ�G���H�W�~���>KW�7WV���cP�������e���\V��4z���&����qbJtG�maz6�i��jS�	h���>]����.ɀ�K���D��3Z:*/%�64��x�=v;$ű����wL����q��xNe�q� -M�O��ѓS��`��A�ĭdzُE8�o!���ｇ�C��@>�%r�'|��*�vv��z˛.>&���Z��h�̀������ߎ�6!' �q��$s-W��h�2�+w�J��pO����}����'Rab(�`���� ���T��: �߯��ן��ћ�J�iO�s��r�hz���Uzb5�� �pP(P�ayʾ��Ʋ�J��e��&[À���� �I�{#�B�~,�	dꝞ�2osS��z	��v���z�J#��:��2���)�c�ع��dA�M;���hUj��#�����K��	!=���r����Zѩa͈�%)1'3Nj�̘�����k����%�3!�;$g4]�(�9��jh�`T�Z? o`J�J�v�:�~�<�9N�
�9���UV�����Ӳ�u��;sū��DS�eɐG�Gk�<����̣@˟�ϻ�p�8�6��|���㦷����ә	�8���⌜T�|{���@�c��2�)] 2 ���ubO"�X7Ϊ�0A���-�UG���v�O���YlZ��������0b_�����BY�sJcC��e<��4�e�ˑ0A�xW����J�RT� ��e�%[H�U�!Rr&�a��-��%�Si\ִ�OZ�*3v��L���qTQ�)��hP�,j�08F�e�.H^�K�sWtf`ґ+���:dްj?�5� ��p�<�*�:\���:E�0z��s�1f\�hv6.�~��_�a)9C7u����tMu�D6}Tu��&�K�ܕ�g?�vB޽���P~�R�!�Ym�ge~�y�|Z�X��2��S�DR�������}|	)@�v�m5�e�y�Ƶn:�ޟ7��_���~��\�6{E�D\z�5u���6d<[��ѐy:�X`��j��(iS:����x�?К�w~z��Y6�F�(��xJz�BO��{��Cz)�����fY	�K�t�Qj�p3�W~UzgK�������+�������J�#����jjc��Y7y���+��v��K�ƸҤ�f9�^8����/|�% n�봆���h�1<G�_wJ�k���W߲��ā@��$���Ԡh�1;MJըv�� �?Y I4��6%�T\��Q��5$�P�4�xo���!�j�(�DQu�<�z�n��5������.�{�䕦�osȯ�K��|�[��6�.�(p����^=�)-�îy��_{���4gN���U!���":���R�AL1�nl��E�Z'��d����|�Z��־�\4���|e���<*Pq����gN<�W�-�Q �'��ji�ki���sl����bo:M�x��I��T@�h�G�X�&��0ٹ0Por6�-��?s�l)�]���������,�p���;�Y�<łW�<���X��b#䔰��Bk��� ����t�)�����2'�";��Q�����᙭=�� ��C4ʢ���mw�"[�������ȡ����ǯ�� r�~�0,lY�5�����g`�I�`��[W*���z t��=8�fSf
+ghxX��R�R��]<�������{>0�A�үg�٭ ��-`��v���f�^`�޴�U�#�?8�§����~slr�"��3Yg|utM��(0��$ȹ{&��d BM��/�����p�P�y���v����<9JK���wI6��DI����AA�B^�׾-��"C���Q�#����`� ?�q�>WDԔ�ȭ��Ź������9Z�r:�$0!�7v��7J�*��;E�%j����߫��3o>����hE���:���ʇ��� �s����n_W�	��M��G�0pڌ#M�&W�Q9�*�uS�A���?��� ~�u�SM�+G�B���*u{}�NPm;�g�B�8��/̥x��)��yN��^=��AoH��L�w�4�+��/��,���J�kr[{7�M��t�X�� �dH�D�|�.qi�}�ot���O���Xb$J���*7���JL�c��*��C ����9��,Ȱ�xcJV�Ū��2?T�-�G�*�G3%�&o�����;�%3��2������.�t����0��d��x_�m��#��jH]OS s�@ި��cY�j��4� ɑ�_�7�Z�쑝�A���>|G��Ȕ�v8V��Ե�G!��
_E�<<#u�e.��5�n������Ā�3��ǜ=�[���Fd��$
��*Zn+�:�j&�����ø-+���U\�q�M@O�F2&ei����]������'���:bcY��پ��:�K\Gϩ{�p�l�qC��l(��WY��o�VA_�}�U1�vU��%�c
�Е�2���	���&��w�Ss����0��ݒ�y�1�V��fY����=N�ɃM�DF1>cy%�c�`b���|XbB�ZƑ�UB"�e�X�����kF�Q����9�GE<�6̅�5�m��������M�<���8%=�z�ɤ�l�L�����ݩ�'�I�}��@�ծ}�韻������������Rc�戱R	�
>��\r�~�0�\��y��G����]�iOt�Aܥ^s�r�����$��d~<�T,=�	�q&���B@���\���ٮ�T�|�nU/F��̕�ǯ����}t
֠��s��D����+�G]k [��/ڤ�P �Y�m����z�]}Uar�1�=r�V��N�s������ nL<^��+O�v&H�g�O�}M �钻�)��D���盤��۪[��o��s�1�x�P O��]����ڌSͧ*����wKc��o�z��}p?�P��-����B���������̬��ܬ�A���,��ޤ�qƑ[
z:M<in��P��SrM��������aK�r�*R}O�ش��8�T�J�袥���L���E�(끕ѝL�x�c�.�5ݝ��^E dy��/��/��Z�# �������"���	D_�����\��v��p��I4H� csO�I#g���E�P�E�����hR�sn��Mc���(������[O�X�[\�ʷn��>�V7���'���7�9
ϼ�g϶���2<F4~���u�0��7��fU�E �O����J�a8R?W�=QU�^��3}AMg��uA�l<xǰ�K��=I�aP���б��[�h�4'��z��J��$���s�/r���ggswS��J�u����Y�7�2��`v-5�P�u^s���{¥���˓
��C�*��� �<��Y���5����0l�h�N���T�9�N$ί�
<����Qx..��b�j�K~U��j��=9<[]t�>�����<A����0E1%�M
�O���f:Tr�fn��ͺ��=J��Q���:R��Q�P�g���m��t��;� �7h7b�5��o�#7�SVqK��$����:Q+�Z�Щg��� E�	�c�tH�X��$�/�&
��x���!�\L��>!{�N���(f�慠8�}{�E$��5��5Ƕ���Fk��p�d��e&��⥹��ذ=�r{�ʜ��WͰ��<��!O�#��ȧ?
�5�;���ys��u��bC<Mug2��R�A\��%#@��i4�ּ:`����I��{�����x	�?v:,P��yRdc-bf�(�1���'�cK�ްĀv�X�HZ*�W��y����l�R!�v|k�Q_ �fjJah����6�e5�l ̻M\)fR��L ��[�����������C~�^�֑�rQym���ȏ�z�3�3%:�������w` B8�y�gI�6�m4�ݙ��:|�9$~��v�y���b�h�Fgk��{��SU�,8���젳vC]�7�}D]=�x���o�9_#΍Ek-2��H�c
X��Ǯ�z��P='�n�y,5噰���"g
���ڲ�d:uώ][G��c�ڑ5��io�Z��9�f 8=�A��J,��N�{��|_�pѹ/Tqt~5�Dz�y_����ށ�;��	��E�
��.�B�F�kc�
�6�S�����Z��P%�ݍ�$5�qt	�i��K|F�S%I��-�W���J��ƚ� ք��"y��4o/�E�}T��[�2�p*ې�P�gǠ۫�K�y���+�ąg�
���]
{-q_2I�̏���1=���J�Qv�O�v�|�����iVY�V�C^yk��\o��
�Z���+�Dv���<ѵhߏf��i-�K�����ŗ�O�\�ZZa��r2���RƠ7:U��X9/����c�*��ڋ���qf'Hjy˝�`�ӛ�	�9 a�i�?(�I�^�iQR�&2�%�e ���y�& �ے�=���`vt�L�_z�Q^ �'����.���y��Y�9	��V��;bŴw���T|�T�G�)�w
+�L6�U7t:E4t��5�}T��n�����#�oC�l��I©|���KK�%�j�'��2A܃n
j��8��S{e��?����c���,B�w���E���d�׻9�-֥ր����v"����T��x��<���N��#6C;"k��CR��iqn7��\��"�୐��<p��C5��4\3&T2/�9%��L*��|����1�߀l�[�w:D,^S����1����Q1�Xy�ֽ<qd�h�q}��~&No�4�����i�g��Z�t�/G&FD��-0S�K��-��!tIb���s�ĩL,Q;i��zE�Q4�'��7K��(ǿ��}�D�;qM �KnP?�R�$*@a��Lw��VcpO���	~F�S��n�,B��8XA'G;z�4C��M�Q�e�k:�+a��3���߾��1-���z�Z<�`e���]��R֛"��ۅ!IV����lɡ[c�#,��oű���)_�����r�ǣld�M*�lG��~���v������c���٘�_>
����h��"��0��.&_�r�>+>*p��Pm���;�d@й?���.�܈ٔ.~�o��}c��ã�Ą�����đF�.y�wU[.&EUٲ�:���a,�����,��{���Pd����s֙���x�(��RQ�=�o�N�L�4�Ԍ�̮&x򣬖@oJ9Ċ�$@�(W�������5Y[T��ǔ?T������fT�@��E�C+F�W��^���8 ����7-I�J���g@���q�ƤP�Ø��0��\v�Dz��L��3��S�я�f"���-�h�z�����Z�_�ʾ%��{6Wƍ��Vv��(���ֽ$G�b����\�Gd�����Ӎx�BL������_|g)��[�)��̎T��lQ
��V�ĕ25:ѝO��+���$�wVtq�o�������$�!�nN^��_y<���<���k��;S���te�"���9�yԓ���) ��4�"�]ȩ���*۰��\�d��m{s�(�!�9��H���#dg�����1��qC��l����@��a.P
{;�t�2OÆ�?�E�k�#�$j�J��+9 ���8|1� 4���Ϫ��P]r�����ypxURE鷦9(�d@���r���`*�yAj�̵M�1wa�����1m��C�����'$+�c��T-4�m�\	R<6�(mq"��L��S�L��zڗ��3uB�F?�a5�z�����Ía�t\[g?y�M������&�����$����.�uzpX��wns��؁�d����+"pk#vژK��ܢ3 �42��)����}\�\*�J�J���@-�}X��*��+ج*Вv��M+@����<%	��b�]�۵}�贚�́�|�i�8�C��_ط����i2/��#b����"��_bo�����k�>��d�G�+bUJ>�N�n�U~g�� �S��7o B�^@#�OO�Di[������
J���qC��7�O���w�ZK�"���NL)Q!�x*����/���@�۠�t&^S��4ė�ʭ���)&����N���H�pO�ns ޶�c"�"�B]K���?0��{kR�	��y:��������^�_�SB��㭗��T�eq��`����WM�/ ��6���D���yzӕ�Y:��-����J�g��N5�8Vn31#bā����'}�xZ|����9MN��5H�n}�$��^�`��b�b�h���:�+��1������.K�����L���g?	'���*N����㐑�J�W��[.V+Ud16,�5�� ;��� ���w_�G4-�׿� h��$B1�P��T��B7�,�M��ߞl���t��3�>����b��c �dZ���[w��x�J���;w��#���V��K*�9p5>i�Nv�)��km�#F����G�B�R���[�ѥ�_y��ͧ<=E�p�#��Ԉg��啤�G�b"�!5�63=�����|��7�*��7|�w�1��`����69>�� �u��
��UnT>��f�Zuc��'v�c6����o@�B�����f��m&�'�	��V�k=P������Г� mfa�� ~E�t�hmq���'/K�!��;�g�Y��j�@5g#�7!7�Lem��T}k8 �L�4�9'�������ed�L� ����ъ�&�����0��c�d��9:*d'Ʀva~v��X�_�M"��	�iӎܚj#����L�G�۾Qs����ŀp_�@��
w�Y^䊷e-�Dõw5��C19j�l�A@��ͼ�
O+ˏ�e�ͺv	��+b��C-����<�۶�iT��mU�<�k���8p	6�`�u貐�D:i�֤bm��`�^��.Ao�M4_��Oz��7.�T8<�1�9y����gx��:`�Uǎis�R��2Gpa��c��5��}[l��T�?`������5'}�V�:��\��'��Sp�4����q4,^���b5SF�r��Ut�,|��N~�V{�7�f����,�����\�zn��	l+ϲdaI�&��:�|`�����n���������!�40���葩+�ō��W�߬�;��*o��s�m&����� �35]��`�E?B�F�f�&�E�\�Ѕڟ�bZI4��_�FA�Ό�)d�+(��uȄ�+_���2�ӷa[j���w�v��-�@V����j��}�FW����?i��JT�-%�n�rY�k�ş�NZ��i����3�?�U #����Ez���� ��y����K������O)�y���:fv��>9�>/j�����Z�(�n'����R�Z֫�3w��:������r+=~U0��lN��s+���#�}�z7~[Cn�*v�2��+����i:E�-K��{p��|�;^�൳��0�/I����������&%�."�����Z�H�L|�f������.QB�[4��������D؆��?�Y�2I\��~�#��YiZZ���8�s�yXϹT�n�T�[�,k�C&�s���Ȼ�> ��+b� !g������S��%�����{dx�)p!tP�:��}����מA2�I�������8L���#�>'+��5�Uu8��*��ݎj���М�8��G��G�R��~8׼��6f�W�\e�z%�X��hXuO��1�!l>���Ǖ�q�7��H@"�V	dX+������A�G�Ȩ��H"��� �V�E:o#�	�|���<�,Yd�pв��Zlp� ��xk�Æ7ͯ�������X���:�Z��o�Kҏ�
ID�������E�pS�y%kMJ�s��� 4y�b6� ���ߔ�ͻc#O3�5ju��0�����$��2��8�X��G@P�a����$���t`�J��|��L~�	�-��ᩝT��#>���2m���/��͐~����-��C�&��I�}��b��/9W%�ކg|�?Չ���ƍ�5CR�S)ާ�RB7BAu����7(�q1��a�`b�&!%o�zP�e��[}��m2e
eVD�A� &k�;��Uڕ!���p��]�����`�G������cS�l��ܹ[?6�J#��p,�4�*�Ab��D����_!��bqf,N���t��9,��`��d����L� �r�N
܊F`<I�Q����.!�; L�tDD~��An�5y�P�5t��O������Y�zn��í��TL��z��!�E�k��?�X�SÓ[à�a��V���.���>I|p��	]LR:1w�݆�����2��ט�f�ML"�4���92�䐥scM��"�q/��1����]&�{�C��ӟ%N�?�����*�1�$�,�����®�!��A* W�S�����wM���4�+�u��)Z֗��AU�oi� z�n�����'xk��]��J7��<���k(%VH�6�$Yt!�
�z]*��
��~,�ZJ����!W���7�~`	�Z�B�����V�cn����M�2�׀���p��Tg_��S���aI]��L8{�B��!ؕ���ϠR�9	�z�9�V�����]0��S9�d�,xt2q]L��!���8�
��	v�Һ
f���� Ԑ���"�WW)9*��Ў�����8R�@'��n�G���>s\���r�*�o�E
��\� �THW;MZ�T�����q�g�{\�������s�����i;8�H�c��6��L�E9�~��),�$heBy����?��#���������/)���8�B�%Z$Ti����X���Ih�	sJbǼ`j�J��������(z�6���w��52G�42�������x�{�/E���;���9�1iQϨm�DKC���n:�u>ߜ��@7��~ ���}���j���θ���=�Z��%
�.\ܮ
)�.�d/|}���QS�Ч�8w��e3�}�ۀ��NPO.�[��kk=��=�\Γ�4��
��]�Sa�$
�S��'�ӸK.X~�`W�nY�Zl�A�#�q�z���kN�ANC��@K�<~]�����ì�m�����ͻr�Kb�1��T��8O�����K�嵳�g��J��./�4��s_Y���J�������B&��5�"J쵤EDص�E"�+�6�����[�EYȼ��h�fH,d��z�ár�����M�t�9l�b[���,�_PZ���BL�)�as/I3|���%��-��œ������p2-A�vG, {�B�jW:�����j�NA�o�D;��s2��qVC��'Y�p�A#��K��DQ=��f�|�ylyL���s֭�E�g�&ɾ��n�`Q��7��������+��Ʀo:l��-�bmX.a�K�9H�zy�Ât¿Vǖ�Ș-�)�J&t}�����yK�2�I��+i�� t/pq����ь9��%}�>X1%VM7]��9�x��ע��H�D3`@/��֬�S&�x*ڲ� E��G�N�F�<��XB5�P�x1vc����J�S✍x	��7cE���P/�Kow,\I��h	$�� �~2oT��
��at=���Q�X��܋�|�F{�tsS�`����M}��F!C�����3LL��= �L�!�(<n����"�V� �����[=�ϲ ���E�\F{d�����ͥ����\��F����]���.���zIϛz:��j.m�a�Ȯ�l�Q6�/�{��U3뢨�x�aΨ��+�~�T�i�,��cq��݆|W=��V3����#�	��?@�F[�g�.6F�Q�1Jn;�Į����_}4��-i�(�ԔMn����#\��Ց�\�y90Y�.���Y�i�pV4���ϸ�4�z�~<�Y'-O���w*��]+���=\W��tz˯�q�T �e\qxcxu.�8!�nE�è��&�9���AҾf�u����G��ߘ�6䀇�A%�r�|��ʠ�[TK�ь~��7m,�[��G���������V,��A��\Dm$3�����S2T]\ۃ*7O8Jx���Y��,I����z��z���<�A	(����9��,��X�J�1x�	���G#��f����9ߧg�5ć��:�x/7��㹐�(vA��xj��O�YcVˑ∽��n��.�7�OР<�Z���1��.spY	~�HǕ�p=y��[g/*����������R��v�1Z0P=A͘k�_u����x�$N,dp�CQs�Ҧ�s����X/_جq�.���@�fh�&�qM���c)9H��NR��$Z�b`<O"�վ�bq�V[dj�����+^��MHU��G{6���~ǃ���s��FD"�_�D����n�M�[Ȥp���\ Aª_˥�Qx�eQ��Y�-�C�*:.�h�8�B 3]gaq�b�G	႖���JI�� �n
wl@�{��JQ;����H��`��ڽ�A���۷�Y
���Z������T�����&����/�)��QS~��J���0k�6(����^k���Ԧ4I�ɞBn�LT��Nu����'q2��Ky�&�f�9��P�xUw��C���i��R�f�Z���^����]�_�C.e���z������V��kHR����S[+$]h�pˋ���L�Z7K��s�@���� [�kA����4�����#O	��;�ٺ�/�'F��� B
�u�G,u�7��Ip��j>�����=�Lڋ38�|�U� �x��1A���y�x�.����a�d�:�8��z�ߴ	��ccb�t���N�(���Mؗ�X���]2π��;.�c�tpЎ7�Q�~9M	�J����"'����	89�bg y�$(����,K]�݊��**�C��ү���zP��o��a����2W%���Z�t.�.����75�0Tx�tW�(ky�$g�4��j�#4�Jw��r��*i��)���b�27��6� �>��Xtg��4v�ݍ`��/�������.�(���v��bF�g��,���e��-d�gt�����P�a��y��p����9�������qP�S/Ө���]
�1P��p4ŧΗp�T�tN4	��u���=�"�Ǒ��g�V<�X�M:�<+�h_w�C�G�,�ԉ޸�POhP�_����e��4j���\��a����H�.P��x�Af���VNp�$'ŭb��&(O�ֆ���u3��֔u$�T��Ab-D%���.�:��}Q�r1\)�O�о;�s�t�k�)"�_����y�]X�[?)��/���5��	EZ5|����;]��F�(E��P�?���ͣd����r��Xx]����{|�Upi7�h},��C����q�~��ɗs���1�� ��G�qz�D
,x>�)-��Ǐ�����\1�E˲g����?a:�U�g�������ǒ�T�3 ǯz����4-�E��C��g펥��N��H]�v�v;�Tl9?�����uW���[/��Wk�:C>�s��2�R?��@�T�A��U�{:�'�70��Lg�y����R\'F��j��w�@fj��
$��վe��0u$�Y�8�p\�x���*L�z����!���ڜN:T~��|j��N����QJj�[��6^'�w���!��:���ٔ���.�>c���E��'C7�b�|Ѡ���[9�j��[?�`	�V�?�|�pP:ٲJ�\TX�SO�h��s����V���G�?	��Jh�����K�'�]���b�PD�t[�<WT&����?�p�TҪ(z���n/*�0��M�{��㈩z��r��څNlNo�ܾ[��|?b�j���I�f��mQp]o���)�-�}���O����7�*{J� %c�7Dw�n�9*~bZZ� sn�/��AIp�hX�Dx�����ޝ&}�Ae)5����%�����g�2���{(&��򨱸��h��?7��;�F�Z�)�T*����kIǀ7��7�v�V}����]:L^�:��WƯ��cJF��܉AA���xg�n8A�嘇�M�#��*�)���pkաA�Pj����Ad��}�2��"��`�r�ӔX�g;v�C D��]��'�I��$�I���G��HS+��?��NZb�2K�ceJt:�o�V4L��%�eԍ����d�9?0�-.Y�����
kJ�
8�KQ��P&��v[��!	���_ʑ�i�9�jC���m�{��7���Jk�눥�p�8�(�U#��_�$����~���êzC�0q�lc0��QÙ�h&�5l��̐,Bt0��a���J�ƽ�HG�D��^K�Q�����Cp��!ez��[،��'"��=�|Φ�; �=�9�K���HA!$,��6E��&�|����֚L���z?�2��nX��+��֓����v\�Ŀ�V�:����hz�,;�5D�iy�/}C�'�/�e��l]����Hg�g�ڣ���ۊ�?�r�`4Ր�(��݁p�Q��Z���	�C��Z+$��y����Oפ1^��[!��>����.�o�͖�� �%ie��>.pr�K�>eO�F��`�G!���
�œ��Mn��!�{�*U�bHO�V=�JT�2u�=`��x����8G���m�z����^Q��k��YN/yf�88�A��q�K���ڢ�ܒU�a����#�ڡ0ql�d�<���|9�E4��_ѹ����Q~cu&&iSZ��/
�#�ԢLY~>�<���{��yWKȠ��؉��<�E��3�g;��m�H��Q?�#lg,��h�@�����m�Y"�N�Awn��i<5�l�"Lt9*�Ϳ�+�!a$���y��V�2�R��Y��>��s�[���_�N.$P�V��߆Ƭp�{P��q��Gme��ئ�ޚ��)=��m7��Mdx��z�C��ҡ8'�����o(8��I�&@n}����&��*�l@?hՊ��"2D�}\�U��Zi� ���Ot�ޞp�̉;.ќ��c$�	6����>�L�����P�|>�� �Ż�6h5�_��ECk+�P*}C|�T�ҧOn�P�q��h$�|����s�|0��ۃ�@�U���Cp�ù6�CoN��WZgh�;�>��s����]����h�ǴY!�~b�kB�0m �4���yj�%-�ϕ��:���![����f�b9�kJ?�h�[�|kd�4�Yf���w*g�N��h*O` s#GS!��9~o���N�Ƃ��➃��?&ޮUa��y�}-�[�L��)���*�A�&aE�-�*|G��h��j�S�yc��5>XW� ��+3@�?(�����GG��u�.��� H���-��g�.X�"'+ꛏi�db���}��F�=�QM�k]l[O� �Y%zdhlHg'���)�n���hM�J,�w�	GL���h���!��/�����r���"�;�H�`v�܅�������9*r}���CA�y�ӫ��:\λ}�A�L�=}~r�(�1�0<k��$�(���϶s�ҷړ���.� '�gK��]��6���0������xL�O<��zD���Њn]0n���,'٬�~����A�;6��U0~{m����T���UjMo ���,0��g��	�g��AtR�]Ս;D��e�t���ע��`��ٱn`ero�֭Sj�'��]G�ګ��a��>�ΓK�	�A��N~ѕi�<h3����%���<�!�G$D��0.��P�;3` ���ѧ���2W�)�5Q���⠟�5��R��[���;�1ī ��!cw?�m��~�T�@�7��Y�kD_w�I�?���[��ٵ?�F�ߨ��'JHm�7�,c�j�����������?�̞�A���?����(�y�|M����u����%0����u�~F�AMg���@#"�H�_�2�&�l�����|r9..6�R,��l�"�{T��_�2㤽��r���B��U\���m�u����g��{p�d�J�#ɨnVΛ����v��;(ϫ���rNY�����9r]��y��0`��D yV���P���ʤ����`��qB��#�Q� � +�^l�We����I�X��B�C;�|���'����|��a0�?�Z9��ή8�ݶڳ.��4f�/� �#٘,�/�7Z�'�Ո�BzmJ�t��
'^���{%4$h7���͊~BZ�CȫQ��>�`6�R6�A�$��8v2n���y�'�r��A�8=��0������0'dj�.pѶ���Q�"�<�2=	i�	(�H����h�D!0 �������$J�D���Q�q��ۚ�V:�"$����IHQ��:�^�>�4F���%m?�%�ʮ׎Y&@�ѣ�!A��(�vfj)�u��#����^.x�]�Q7�xQe�Q�
q���͢7Q��v�M�P�kL�'�������:��&Q�,�d�ԫ#<J2pK]���l"� tg\o�3?��(���sd����/���� P,��j�<��r�>a1�ZBS�#8XwV�����p���#K9�Q@aBxj����'9�
�^B[؝˷<�5Qd�&!"�r��Yc��U���S0�Ҷi
ͤN��������ӧ��=��g�V�ُ�Y����Q�y�kr1�z�(����&	����m���SQ����ZDh�PU��	بӕoF�BwC@Fן���ST,n�9���bBB�o*MlݨR��6��0�����3;m�D@�Hܞ��`�0��K)����r��Qu)�zT�(��e]Jwxj+Ғ�L �ܙ5��ӯY�w1?~�׮Bw�!�Te�.��,)�����Q=04���T�cc�����l@��nz�dʅ*�јIh���?�]Hn2ˮ�:�����)�\��fo�_Q)A6"KK�3���3�=�Tg�N�xowi���_	� ��n���0�b[e�����G�׸�2�e�>�_�x��T�QV�� }>1�Z5?9�$���UG��o5��@.?���K*ZCiR_�%qD�!�p'��ˏj^�:�=^X�W��R�hD�n�&1-�G51s��7���{�{�$���ӻ��ϒp�<��b��ĨF��c�<z6��RY��(�kfR7֮��䅠�����htʌN�٭[1OY\h�B�Ʀ1(� vs�ZO<[\/�YxxL<�#k� _��u�[�"a��]ұ6�p���U��g��ց��-�k��bel����^1G��G���T&�%�#��R�D��vIK�������~e�>F�w( Z�+:Wz�F
�dz� �֊�j~f~ey�@׀O�M�rT����<L�,�5Z��Z��ց}E�ے0%k�_�U1����N6�Rb����V^%�̀[�[�'{Ii7|,�K�W)h&�	�����X�G��ɧ�p������c�&8��/3���#]�U�B�a2�� {���h��:�\�z 2G8@y8g�������q��2D��q!��"���(��,��-����ؽg
2-/��	^^p�L��Z&E�x�� ,��\e�\�9�Ck#~Ea=*���A�N�O���I�Kjq2t�r���Yu�&�/��T�S��S^��$;��V���aP��ےlS3�Y�+�^J�5'A5g�!*�ӳ�T���϶����揲b��R�Q���q0f�5e���3�i
��+H=��/�m@+A`<�m��ǋu������`}��� �n^tG�e1d�|�\1��}�́2�_A������V$I:=���\�j'�iG�!I{<������|�r���L�N���h��Fm%B,Ѕ��n��5���B��M�=R*��eW ?�0�U���*I/d��'/�����
,<�;��C�kFa\����o$�+���b���x�~x����q2���[Ą��ӻ��_�6�4T�zY�Ә��4G�Z����J^�H�UI�Y�w�H�v��w��r$�	T.�s,��4����[d�a��)ʁ��N#> �4�A'�Fw��N1��yO3��Zf���f�\�_�H�Z�a�
+^ë��9?G%.�8#�#tJ��{{��*����u���C�KVZ/�K�*�(��,*����i��JL�������ɐ���C��ɸ��V�1L�G��д��_3+��a'*��o�����I"�/��.���.�Rm�hc�	�ɊK�&Ax,�QP\�~y��ض��� �VC�Q�U���r�9G��
���+�**�'b��Ҧ�WuX( g����t�e|3[cT` /���h�X����؟ZE7=I
\��T�6+�%W������iP�p..�  �/�
���}��{�B��a_u�}+�8��`�@Zy�oCc��a�(��0�˦/��p�3�o�%�0�F�f%RQ�3���?��p�5���Q��d&K��.���g��="�TD��\�R�p��6dE9�W$Y-�x�Ml�r���VBoў���⚖H�r�嗃{�P��j�^F�(��s�0�W���^R������R�F�y�y�}95����cF#�:8!8洸N.!�b7�L�J㕃c\�-�_��i�#Pٵj��PX�����m�xv%�Q8l%N|����E	�iwu�QsS6C ���C��U�w��NlFP1���%�ٺ��PS����o��[���y�ގ�6�����v}�ƻ�h:�>WO��Sޕ�����[�=�l�!��D�AU׏�G`���0�ǽ���9ҭUQ,G]���A�Z���bc��dĳO9�J��}�����F?*\�Ȕ�LQ���яz���J�E^xF��do��*��FK��N�J&A��dL5�|��t��8V��u(�������C�AΑz<�?�h�Xs��;[��M'h�A�o/.&rI4a�E�T���1�@��Qdv�s�����DVBp� �53sehA��F}Sp^��;��a��}{Y�u�;��"׀G�4E�ЋN�ލ�k�Y}o��J
�@a)�)B"*Z!P�%�F,�"N4�W��%�n6Kg�șѶ 1�b����a�x��	��S�D'�:�Bn��_�Ë|(>�\<�jLp���-�?X�O�;4V��b.5�"<�&*������G\.>h��"�^*�[ʡ:�^w�/ �e�����.��w
=6��k�Q%ȧ�a/���lD��ѿj�q7�u���f�[kN�)]G��~~�hә'���p�;X�m�JX ����E�5Ǔi�xmus�����#�UɈ��zt�9��N�r�ݎ_9;�ڎ�c�V;JWܣWW:�-�#BL!r�8IC!L�O�X�<�����<�xJj�ⶦS��@�ZL�j�fB�2)l��@�	�k��l�9?uFn�>���t�S��a���--���<�Ť�u���J�Q7�n�	}Q^z5f[&�M�ٕ���T���,5�Vx��{(E#�M�≈�8�|ѻ��m���=mt����xF�����$�De�!�G8)�9Dx֦��2%r��7R_{~�>}ZSiNE��ެs2��]��۠1�}{��L<��^�����|hX� ����m8_��ȳ�I�J+Ϋ�&�8vל���y�(��K&a�"J�
L%�z�߬�*���1Ȕ�<(�}.����.I���8�C���Ò8�u�˨л�ay`�za�-��>y �4�Ǻ'"���ʻ��R�sD_�f�Xs�h0(wV�A���
�,���ӿ`�m��Co��w�{C�a_B���*$2%�j�p4������%ד���7)d��i������J����	��*�gq?��b�Hy�Q�bY���
�sqZ�=j��S��bѵ��r�� 'A0R�;��JyK$a�P��J�*k�r��*��t�==��ѝ� ��	�fpSqx��dE����!28Z��y�tL�M�)��S�
2���w_�w�Q����0�u<�n�;���� E��>����#X=����Er�y�[���m�����Q%�M2��{�BD=��ʧK>G$,rW�W>P&�QH�ms���Z�9��t�~6��:lO��t�tj���M�c��;
*Q�����¨;�ѐ0��s>X�GQ�1ù�T�ÒI�@	��I~k�^�k�J9y �nK����5�|B�¦���2p�8��~w��[�l����ēۼQbC���K�]�AËb��\��	-�a|�5�ߏ:@�$�.!f����"9�!����5�sp�z	^e��ߝ��GIv)��I���U�ۄ>���pZ���,��d�g���Y*M&�$�	�M9�er��~=�U0d����4?�0��`[Z�	�v����٠����]c�ӕ�v�, ��]������z�o��UxN@N��X'��P�81�_��^�.������*�U����&f�*{_���k6@�[�.&�싇w��&������F1\��b�9�K4h��r�U~���m����.d���98�@�p��lh�L�
:��Tj�!U)8���#�y�^+.��P1��]��i�8���SA>�6`'����x^�t���`c]ﰀ���pn*��k6�Hg9�G����[&� �[���X��7��� $6LN�ff�|_@�u��W_	��U�����E�:sBh1{"2:��m�H?O��%���U�,B��۶z9�(Ղ&w��2�Cu���R8Ly+Z��Oa2�"E�)�^怹�a��ߕ-�!QM��ʔy����Z��2�'��|+�H�:=NǪL��fKA<�~BNʤJ��{|&h����@b�)���M�G 9�"��+�W5AI���45��k���q�4b� �Yq����Qv�yf��I��L@��*��/����C���Hz��Lm�Y����gOa�^,��qP$3�wiR�?�Q��w2XZb�?�V�,�?AUl�xT
���	�J�7W�y3\��=B�D�V��R���T?<@w�&:ʦ�����?qa��tL�Vz(]��w���/[.�X��w矜K��Ad��`�?�+:=s8�w�&�&-�9���L������������UB+�������c��MQ=�4��j�wDe_��G��@K�8/��hj�䓄(�����!&.�4}<w�=��H��T�}]����:�Nw���lg ��+��[M��e��龦q�rg>q��G=}�Yݝ�k�O_h��r`�������$�lCo{��n���j
W8��AP5h�:]���M��X���lLd�Q���� 1+)�	��rV.�n��*�`�rS�Hǽ�&J��}�ύ�G�ݲF�����p���"�A$YS
�7L��&�w�/���{�Em-[�a����c��֠W�F�ڏ��Dsi��8��;�SI~^��2��=��w��н>�2��
8�|~%%*�*�9��h(	�0A��h8�"H���KyT���z����������
:�]�$�4��<s1m?�h���DS�Բ
� q��)��?t�
Y�㹒��}<�M�@F(aڙ)�X΅�[�ϙ�����4A��R�yU݈^	��lJB0�$ a����]�W4K�f7�i�(�;`9�ۗ�[S]�b��yr�3���z��#u\����{B���̋�"J�YK��q�~��b3�x�L��ʶt!Q�S�#+A���4�pD����6"�w�+��,���-�l
�g�\}V�u%����/�����H`�j�m[M]��"G9�:��&��1�.a��$��A &�&Id��w�7p
���9g畬�۱o�������%p6��=Ǟ����G�뽼r�7���<
%����Ŝ{��u�\��T�2ĚA�l�О	[em®��V�/�I�_.�_�����O鸒�u��b%�?��S^e5��/�����^nҬ�kj �VT��r���޲����|�#"��U�8^�M�fDN�-15w�~��:�ˎ4ǜ�z�a��V=舤�X�ͽ\�ƹP0����w��n,^���qD��ϓ�H2}̗K-J�n��z��N0M�
�S���.9*���B��x�M�"�|.qH��<�Dō�ؕ���iK\Q������m5ܮ�5���{ ��^�>��|��E!�W;*h.D��WxN>����Y��-�l���׍�������yJr�(���jenrto��V;�whE�4*�堞�Ĺ>��3mAn�K�_� 7��d��L�B���(��i��S%�^�ɥb�XU�1}5�r�_����޺��Jc�4��cE��c�f"�5�b�yǘ p�I��+-�r�ޱ�ٷr��FS8~j��G��� Ԋ�a��� j}Up�����>������ �g�����8a��A���QeI:���C�^C5�D��iv��
����=Pm� Bu����1����țeb+���YE��6����,GF�Y���8�q��ԥsL])w�ձ�����C36���d�&p���uukg��ѓ��x�r�	�ա:g{Ԥp*�@�)�=S?D���c�<d@M���c������,ص�e���z��r.$��̻���EnD�Kp�p����m"�{X8Ur�$�_v�s�r�m�Œ��P(0�� �Ҏ�������z͏h����ZB~a�r����߾��b����m��gHm�fo5��W�fEQ�A���C��k��u� �Ð�<E;Zvl�d&	�T��$a9���C�"�)�Vqvyf���1��\y�&@� $��Rԕ[�R��n�~ �$���b��S���y\���P@[�(]�$^�*�J�Yo��Xw߾s�e�d=���$��4(6�ݵ.D �ᕃwu߼'�J�7�%g�Fۃ�@��E�a�'W�0��i`���J������H�X���>��w���K*��
����D'sYZ�bx�i�zc�n�w�I�#7���HQ�o��; ����&A��%`wŁQ^)�l�f�b���O�>�vp��&�C�7YI����l̈,�E��H�9��`��.�p���B����Og��9�ˣ7��V�J7�6��K�F������{��6ɩh�h'��(�#9Ci�w�J&�J|�4��֫��2恾瓪��M�	�4��6�diI�������&���yK8����'��Ӝ{��4F���qoɚ�-�Z�:ܝ�3_z|Z�L\���h�c�L�+�Ц��R�l��ܤ`$n5߽�T��0���F��A̐\T��
T��H���H[Q��F�F���b�N;�+x-���=�n2+�'_fV�c��`�]K��Hӄ�VI�6�b�����Z����EK��V�$暝٭gR�����@��H���[��x�Wmi6o�Ku4R�w"3��B��c%_i�W��2S�DG��N�����v�G�gL]��8���t������˷HWp�*��9�ˀT�,*و����jK�0obo��R�3�)܉(�Kq�W�(�P��^�XC��g���C:Dُ��@��s�|��%��߼�1��*�WUy5��Ř�.�C0�@�lm��V��
�I�o���ó+Y��ޠ��m9w\���ҸS�T���Y�i�A�*p�%�C>J��v�ݓ*�	_�N;{Q�r���#�D���������ލ(�c�{��)��-���'�ᤶ�E�y޵8�����ȡ���{J��dh�z�&�/��Vt�!n\���զ�򥽚se�:���.޶oBcnHQ�~�?�}:b��d_K,��|�&�x���+���4d� 1�����=9:')�`��z����<>Gy$�	~��}�J�G��A����/�P0�(���27�"�^e�
�0��=땪/̰7C��^�"¬�eG�>w@��o��/�c�=є��M\7�m�6��s
b��rn��hi�/�c����ֻ0�"����h���@��n��c��9�īZ�̽F�O��곆z���N����O���Q�'UK$��s;l�U�+�
\���\�� }��)�Ҧqo3$������{�Fu�ӟ��]c��w��z]��bԌ��im��_���z��� a\�|l��� qjN�0� ���������x�H=���ˠ���Ea�3=�G�)�d��>�9;�x�JaW��{���fi��LPI���t,��^����B��������s��&pa`=t���UZ�	�M��"�nz������{�ꇏ�Z��w�5�բo���uϖ���72%���m�&���W�B�K�%�@z��T�b[-؂�>���-��U\��b�k*��Fq���lУ�Cn����2W��+�
�=���
��~��aA�O�iDTUQ0q�nd���m�
g�*j(]�x�+�2�Y�lȒ�����=U�q�;qgȚO�ؑ����b���B�����g�( ��ȦEl*z�^<�ª|�cх��|��l��3�L1�@Ϋ��C8[c����嗄E<_�rW�B^A���<-iՌ���Tv��iK�?Ş��305I��(�.(�v�Ҡ�LIqԄE�	�<
 `���{nox�뉨C��!��͎�����~��{���J�
�;�����>���2z	����f-�իC��)"kmǶ/*0ՙ��ۀ�E�Z��I�,�SJٵK*�
��]�5�w�\&��v�Ҳn��g��am���8��W#����i�:ީ��<�S�a�yo�
���\&�Qku�?��a�&
���U�a%Y�21J��p������&�n�I?��ݣ>�AZAl4+�C�ܡOt�����
�"A4�7$�g2{˞�y���ă���&�?Y����}+fQŵ���~@Ro���I�� G� I���*�<��#�Po�lt�:�L�L�����1����~�K�Zk����o��vs~@���[ 6���`�#J aXԪs��4���P���\^�,�]�z�.>�vX�� �F�]S��֧�J�E�?ܞ*J����E�����M����<���A���i	�#�1me�H�����%F���l�o��YUg2���$�kz3Z�r�J)K���V�\:��A�[�F���i��l�_M�$��@��Z��N���'���M����j�B�� ��SÃ�k4%[D�|$Cwo�X���(Jb0q-}*-X{e��ғ��+$&�V���bV3���F�4FS[0P̞�|P� �6��B���ʷ���d@KQ �Lm�gB����O���@4�٬�Y|9Y�5plVJ]��m�	c\_M���~c����{��D8e	�YK@��
����t��t��Ђ:�6`J��h�B��f��$3^a=dz�!��G\4��-!S�Z�,���ff��m���#��b�K�B̽;��Rv��B-n u/�K��]�Zl��Ȯ�z����i�p��Z��]�*9b4>e�ю�^���[��|���y�'Gۊ����O�<��z"���:S��[8XO�և�5����xg�����&���q��'�H�,5N�����*�bd�;����y`�d��sݯ��Ź[�����T���
�H��ou�Qr���rn
�	r
^�����4ztQ�Q{��hl!��@��X��:��rE��75��J�i��,�=[�}fW�rE����$�zrsB�io��^���wE���=��`$+QK���S$����r�U�]ٜ0���5g7ӳ93�$���F^۞SE��Qj�j�u(&����k����㪕DVb|�R�3y�Q��B��?�s�dUy�5A���g��čA���������I��ԯ��n��d�����N�/�p�=�$+/�F̛��"�>ѝs�ɘc ��o�s�u���P��ݛ#Y����37����v�]�J}���w��3�qej�!M.v�b����%��27jv��ɿ���)�KT�����h lS�X]��-3�#I��Xp��ʴ_!��
"� C�m�F������r�w�E�c/�=��;�
��&��B�ll��+�Zկ�C�t�+�.���S�iZ���g���`](�G�_�� m{�������a��r/��AO5:|چv:��z�M�xgaYjg-���$E��GX�V~�x8PMBV�֜�}��b���\�����z�B9R	>�+B�?h\io9�a6�[����iœ�$�Gi  	r�S��E{V��a��m�޳��G"r�,t�dl����� VŗS���
�Q�P���pr}`��FSu\L�(0� g���#?/���*&3��\��yP`���9�Fl�G92�:���ӗ���1�]�^��:y�x+B ��Fj���� �������7����!r��rk���W�C�W{�k����S������۔�+���ش�)$�s/�Ks�v[�V����}�H���u��˶kO\�1w��E�/mP8[{5jEw�qA�<f�4iY9Dl�K�	�� �K@��nJ@���4�l�d�#�E+�hs�Jm�ҫ����������{��<S�j/�Ɩ8D�i/��UN(�:4F%2���Z!K.a�q���{H.f3YEoN<@+��\I�"�\���<�Ee�g��ӊ�b�8~2erH
���AꖽH�,�V��2��}u��7;gy1�9_�La1���Pn�u�%ovƨ�v/�m�lff*@巌N!��v�I�5 �?��i�z]h��K/_�iL9����-D�ow�W���N�����?#�,�@��Hέ��Ǝ�"Q���>m;_��f������O�X�V��_���@� ��
[�|S9�$4�yͼ�������"2���3fNF�&��0V�G�ɔ$���<8�F=3�E�GCCD���	�lU0	�+��p�����)�ɑ�3��(����c�*
"-W;�����.�'r��!��	�JA��ĕDώ���d�(���x/�y۴sq��'���^�����
���{w�8�r��%cw���U��er�!�В�ծ@�?M�׉8�����`���B~�X��~�4�ӑx:��q�ոo_�	�����b�_�uo�3��	#(���k8��q����D�Ma>��M|�<��f�A��G��S���]���a-J�좦5�#:f�)K�}�_�����g��Fyr���Q��0�hrN��7uw�6��_19�󻺖�&�b�+�QV���-Zz@Q`���Xퟨ�u3M��H:��/���ŉ�����ldr*�` aA2���O���5��N<��q�:JQ"�L�h���s�Y�$J�w�G�y�rJ̹����Jc;h�JdT�[�������V��2��y���H1ܠ؀Y�E��C���:�vf�����	����lG�Q2ӓ���E-�1�q}���Q�B'?7�i�N��TX�ԑ�����~��L�1�"�R���r�q���+t�QCW�d��T��p	=��!���:�#�p':�����۽ti���,�/ �8$����+��OE�9�ɏ���c�bTC��)�t<n訩C�|S�Ū9[��������g~��ZZ��P[��V��,D -|x3��$��g��ƍ@�H�lD��� ���z#�
�&6�!�U�军=	�b�Bi���#���y�@YK�>����u�����*�L����]pK>� H�6�P^�R�O$T&E���9wQ}rW�r����WH�)Us��V��2�=�3�8n�+���6#O�/_���&3�AKc�ǈ��|C��ji�;�s�� ��
�ЃW����z���Cu����$��n�\Bìd�P|�d��R��FÊ�hs�tHy㵝��[(��-���uOַ.6��?�W���-�ko,�����Nv��#��o�51e�����{G�Id�*,P���sM���J8�!����R[� i��3N\EsiW��:�63x_x���ff��fWV�{C|��*>>#;�}�Ȼ��9��3�JXmߵ��>2`���u �^_j��`6�e��x)�٭��p�J?]Z���.*F�*��C�iT�˗s���a�3权��::�]Ĭ�F�!���C���}�����3.����~�/�y�q�� $�toQ{d���JMW�3W����A3���B�u-0�2N�0�pEA'V׊���a�pK*�>�h��2L�Y��+ '�s�b(�D���[����"6HL�om@w����(\�,�|NAL�z�q[i�E�{���V҆�.M�O�v���a@&7:_�;a~6�엝[�19���V>��K���`�ۓ��<��LCm:`��6�"��:������E��z���ǲ6�l"W�Y�̨&z���8R+-<CO���L�oUG$��n8�ѭW��m��Q5����1�b&����Ub�GJ�X�'�_��UsΜ���Ȥk��&3ű~i��{��B�\۩�Dh�~3�)3��AdW���'S����Y&:=�lF��^,���$Ţ�/��qL�*U;^Ӆ���zd�xp��ymI�V�r������Ⱥ�H��y��[����d$x�[�I%���55Y�a�ָ��p���CW����`6�@�39'��rO��
m��������R5%�*��`V�� י���R��\@[&>���]!���Ͱ��n�k�B�O������p�JI�� ��hofW�I��t�i��)�ҥy�t��3�h1��,7�<�V�1N���p� ]L�mnEI�F��PR/���N3�>��/(|�n������bM����L|�*����g@8VV<׎�M����|�<��섺��~0�3�60c�E����O��)$��pʭ�#��u�Oc�a����b�Q�`L�_Q��A��,x@�/�EbTZ��z��Xb��T��Ym���̲X�f�^���J9�tJ���E�ݴ{j�Y��QU�_�fU�Rru����e�Ml]�wo�>��r�l�.�p=�;��?�j��Ej[P�;f*$;Оώ3(�SYTg�~�I N�覹v�a�[j�g�"�]\,�r�1@C���؝�bh`�*����?b2��h1zt�9����?iO��	�2ɸ�Ao>���M�xp|��b}�_��e�;����ă�m�;�3 j<�r���ǯMd���l2?����u~���G!�ȗ��0�^.P���i�� ��ʁv��Q�]��P�ت;i��<�G��6eG,�18��qL��Ur��[��?�J��)������r����ys/��Ph��]��d�D��4S:Ӓ�Ã�tz:�y\7��6�|	'X���9(vo�mi�k�\��	M!��Nꜭ��2�T>�0��|�(#q�#"�'3&��0ȴB��X����t�qK0�~)1�u�E�B���}\�W���;�O��a��oT��S,$�#r��~�)���qV�㗎�R�.�Q�����^�VHP_�?���]/_����nQ�48s����5�� ��e8�&�%f/�<���٠_�{X�HM˷H�=JǪ��L��-<�w���hҹt��s��ؾ�h4p�m�����|�����h0OfA/���,��`*��Ʀ�"� W��EJ�t6 =C�'���fwJIp�M)02<���t�t(��(�l��jie���<�N��|��F�<�����ʒ�k2{���*T�~�銎P@�"I�A���L@�����M�?��ȫ�R� /��y����hL	����T�t-�'i���w|�� ���ퟡq�̓��~����71d��CA����%��'�lw -��/�����b���$E�/\O�T��$���@� ����]I�P}p!@�����T��X�v��/B:���	Q#���m�A���$	��}ŗ[`��������l�L���^h�W���$���a.�ǖ�z�TT�?�Pc�����QC�A�9|U�-�.�f��S0���I_� 浽5�щbK3I���B_�ܾ������秉툐��.I~~/4�ɕFd�|�x��% �]ʄEu*/��4�6�oytY'j\�,m�h1X�����8� E)������xѯ��f%�oC-����A2L����.ƛ/��˒�tt��ٜ�IQ����0����Jd��3��0óT����j�y`&M������6��?Ge<y�bڣo�B#��_~$vϻĬ���G�TT�]Y��*V�$w�k`ֆF��6/@�U�-����'���"��^��}xy���g�_a Fg�iJ�ڒ�����"##�f�����gH��n�8�za�*�J�d��z	.�ůFbI�=��QE0y|n�[��n��h��K�R�=C���d�:�`�D�狦Ux�R�F�B�#"��;�w���	���V�Qk>5�4tf�qu��-�����lxM~����cڈV�����J:]�4]����\w�b��T�?�v��%�ž*�4V�}k�,t���J�	����5���k��AD��冚��߄�ҕD��X=����j�0�9���{G�W�)^�"Q9Y��y{n��*L>���1a�IՋX��+�3�*�/�J�<s���������jL�
Pw��c�D�5쬌u�{%�r��m���>�^)m��e<���]���uf�L4g� n��H�$���e�=���O#���������M=$!�l���DO!=\�k��V`�̒HJ�@x"�\Hu��b��3��JV�ԡ�a�c��%�;�wl��,�R���z��9��U�)�o�ױ@.�<�V$ &};	wJ���J��+I[�(w� �~���(mc�N^���P��ѷ��Py�QU�����
���=�^��<���Kc��y����ؖLeJ�=\{Sx����N�� ��k%��>C��A�_�hԴ�._��~+^��J��u�~D1s@e~�LU
x	*"�Fr�h�i�D��g$�aB�{)��{[x���Y���z��R��+�]�d�[�.=�cu��yZ�#�5���G p�g�[�G�����CDl4�xPb�G��+��md@��@Κ��\�1���G#�]�[�Ֆ�!�{��d�A�J���1���M��W���z���!�^��W)I�4��9e��U����8�@CI���D*���W��a���K:��GlOIz�Q����U�n�c� K�5*/�8�y ����ȝc�O�B��Pl(R}i��e��!4R^��f����C�9o�l��J4(��{]OI�8 ����?} H(�����җ�g�/�%�ݴꨍ�����c�c�b�/#��G�&�!k�(�V0���-���v����RN���ҥސ%��S+;I~�_D~z���(S���ɚԴ�ܕk��#W؍��DJ�� ��.U�Pޙ�܏��N��v�a, �8pȼ�V�cg�M���DG���܄�%l���'�O_�)X���
�jh�}6]���ۨC��R�'o�������f%����JDcDx�y������g�I�3�/pz�6�n�������,��9OE�ϴ�����W��b���~�k~�x2����s�-�mQ�=����u�(�y�D�}��J�j �[�6�ĜU%(A�n�:�R�>��v�@�oDK�b>W#˖{�x�X<i&KH$V�G$�9�v�pk����:��~�m$WQh�F���������6�`A�~3�+�GOF �t�s\�y^MUwޡ�W/
8̰ =9*��82��]��^��������\z�� *�����1��H���`Y�Q�a��7F�4�2�1?0��t0��^~$�n�L���C�]=}�T�Z��7�g���2�/⾗��A���;<O�G-��a�J��6д��!�O\��p���~���
9p,�M�(���]8�j��$�>�)V�2m��ҁ��~yRDE�$V�!2x�&�.F�Y��z�%����&o�4����a7ϻKN1�,�n��w��?��?�M
uΛ�,�����2{R���*�hX�;���F$��W%^u5e���M[k��vQ��L�f��Q��m5�'�`o���Ê|�1j�sV�I���������2�B �9��>�+����%�',\��CF��a��	�hLo]�T*�rz�6N��*&n������"d�ײg���	1r�4iyC��;�AD1�#�f��iX0cb��q�N��6�s��r$�'^{�p[�坁�� � �~-����t���@��ѧ�sc�_S��T��#¼�5l2<��)����'h$$]�J��b����zY�w�*k9YS�	]�c�\Ac����%�#В��s�e��Q^�����?m.pr���L���^�����F�e�e
��	����W���lA�,)�q�`�E%�C��A^iB"��u`!҃zc!T���쉐?�1��'ߛ(iM��m�
h$C�O�� �<�b�w����WY:|��g�H��VM�2���PZ"i�b0|������m`��fFB����B����F�F
��j��Q��+�NeC��w�~�1�I@s��1x�`�^#��2FmQ����뙓�5��ۓR�L��TR����T'�f��7�$��}v��X�"Ll	jx��JE!�r=��X�ޕq�XuOG5N�}T��cJ�#�B�N�<��["[��Ka�PB	`��=�Ϡ�N�N��04����܍�dA��<U�Em�l�C��$��؄��eߡZ�Ӌ��.��ɾ�u+o� &V�Y~�<�q�}��
��v�/��5���Gu1�A����a`����D�0M��]L��p�M<�	����t�{��8�I�>���x BU�μ�f���.UꘚL�ԱP(��b����Lp�u�h�|Џ	o��_��0��Z�]1����2-��"W�^�6+�h)_5#����E�1�ޑmp��L@-j��5�"�j�d&��f컺5�27'1�^"G��L6c����/�$��yy?������@���\&�v܋cw��P���(N'������{����݇����0Taez1l���N��Km�V<��/MS�p���q�`c�hRN�6�����EL�g��&
���]�&[��\���}V�o���ֈWy(�tM�Tx���A�:�x߮_�3����$l� +�zO���h
�����og�a3P��q�D���˷���)����-�N��R���}@��]�>������k��6"�.qV*���F���RtAh(nS'��v${]���n�b݊�{5 ��tO/J�v0�M�E��7��Dg6��Ǽ�=Č�'Ħ��@rt�n�e�;[�*��>ܝ�_��l$f}�+w,�T�R���f1ꓱ������Λ>���w��b+�}~I�JAQ$x�I�һR�0��].��+�����A�YE։�(�d$�\�hî�;�p�F����ژ&g��_8/�~�4�h� ��Zӗ��VH�(ZtIT���`��@tq������ک�ҩ;Pe��{đ��x���'ƟF���I|m��O�i�@��p���oȃJ%���J&>�^���u��d�,���3�qA�JE@�}j��y
p`A�VTl�X���DV,�Q���X���H�~�Y/�� ��f�h��3�4�5pZ3Z�]kC�?EEEx��m���6(mߏIC��5����ɡj�X�b���������w�`bͩv�$�*�8}2 _Б�FVl��aU�Xc��E�k�S7��m��j�z�x9��r�_w\-��U�)�k;���/��1E-����B����X4�71�K��ysH�}f޿�0����&���e����ŷ{M������78Ljڽ����GQ��L����\�I?������ ~�����l�MZ4�`-��!����������vاF��G����Q9퉊������h(A����?*�ҟ�'�:�7��ς!�ڝB+��m�l���@� �Z��t�P�Α�Βv&�3|.D�����V]SWV��I$ۜTC��Z��^��
8�ƌ������ ,�%3i7m$H^��Yl1X�r�3dp�U��Cء%-d�]�pw��ޢ��@�UK��ů��J�c։��+�* ���I6fI`	��nd?R��)=S�_{W8�e����k.-����ڇ�ҭ�e��A��$���F��w��O3׿x�`^sM���`��{������b�f��v�ǵX!��O���#$�Z�I#��{���В�/�-S�V���Y�*��-�&wN��.6�()�;��#�^>T��p��3���Y��~�/hu��SA/��;�xC����ׂ��?}BV��v��t��T�l[`��4���hb�Te��Ǎ�tIw����^Җ.�����/bC6���Je�oo]�kz��\m���Z�<]h��<D��\��W�J��!��1�o���"��6�2��єP)��/amT�˘n?��D8�y��= ���9�t��w����Yy����;E$L��V�[l�~�PRQ������Ӛ�����f���G���lڭ�sԜ���	�����dJ&��k:�m�6���|����ܵ�־�
)
՛�x#_l�v[�\怶^E�F��&���>�^b6��DZz˹H}=t<��&�ު�>��v�`���.@e�(]�GC6��mW�ut�3٘�����`#����Ak���L*𯅯��cΫ�����`���íx"yi8��P4�QӮ��݌�ã����!���¿�m[↠:�Y�s�v��`��g�A�?�h��a��<~:�\o�Rj�y�fve�@IP�tb11 ꐎN+̄X3sD�y��9Mn�m��x���-��vi��L\��u$�u^s�<�c:I���{���L�c���BH�\|!,�W�"$���˅���`��7�) bQ !��x�B�촻׏�(qĎ	$͋nI��F�����ϩ��Kz��5ꎣ(��z��l�H�Oq��N�ô����oPI���hTԄ�Y�I-�:���g�5������='+�����-�r�v�{-��G��k��D�{���G_��0_w3��h�-</�P���Ţ��mm�ܨ�>5�^�����`����q�|��17i����F3�w!_@����ь�2e�4��}�)|��K��-�c����e񽴫"_U���+�~5�LŒC3r"ղm)͂��Gˊ�K��G�qH)A��]$��Nϣ�)�¾e#��������1n,U"��{�>{�.=B|M )�#?��.S��OI��=@j���J0�)��PU��x*��Z a+�dS���Ų�R�k�8z��P{}b�*sQ��S*�3�Z�]�t������ :b7�I��B��A?����cA����p��� 8��F晅��u3���ZW=���	 �R�b@�X���oH`H����q���w�Y�b|����lէT�Vr��	R�����(v�jA�&���r�٥�����N����)"X���A�w����~�����_%��޼U�d;��C+Ǫx���;�nhq��+��[�\e��:r.���@�y=)y�׊_��# XiI��ZD��|he~�l���s:Ť"��%8�z�٣�T���N�צ)J�v��2I���p�;P��1�um�V:+*��!�4��j�V�����@�0�"���-�������X.t;~�Trᅱ�U�O1M�66�+
|��*H�����`��}|�=8)1	���4W ��f��N%f'�qc�2o�{3raQig�&9�;���+�z�/�gJ�����K�ca�$w,��84 �L��?銓,�w�f`��
�qbK����īUTY�@�l_ψ���Pv�ă��0�N}᠜�i�3"c@V�<]��ⴎ�~Og���_�P��`�� 6��d��~s�
iۓZI��op�앨ts�Q�EH�N��U�ֳ�!�$��j�")-fOV�9�����)<�1�έ.i��}��T
�fNG�s�7m���P����9'�j0�mI��O}s���.0?y��c����M�4`Kx�A�}i�N��i�����_o1�7"ͬ7�(�4�Nb�\]_y��އ�nơwȱ�|�&`?J��$� �uAJ�iٴ+�y�TK��|6q��Q�~�M�u��^J�{�A&ە`9�d���"�� ��/a��c��4�A�
��y��h��:`�3V�A��+��=Ro����vO���&Y��󟤣�^6�>G���RE Scv�i����.;��t[��,cV^�~�_�i/t���f��·�g:��nm��%tB�[&��#!�f���[��<�!�FZT5��!�/�+~o?�mڇ^�`�a�m:a�P���c)�����n�^�g*�V牰�
6�a�i�p%��  C?�X��p�]��@�B993ka[
�S�@��l��E�J�W�`�J����1��&&��/금N1*���Tz�kY�M�?�E�(]�;�G <iݛ`���:�)���2qa�J�'�����RЄ�E?��!��Y`�� ײ��
j,��ƶ�%@U��A�����;�-���;T���m�*���D�H2�g� �D�=+�aNJ�6��6�jp��@'~9���~���|HZ]5?��hzW��3��E~!�����Jh��#��O���(����!��a�Ƥ�B፭�����NVfI��A�R�<�D8���!/��c��2
H?�ۨ.Ё�ↀ­��#6��!��jD�S"��eIǱ,_�G6���fΑ��&���7p�Fn[xގ�HG:M��K��;h��k�H�ޥ������
�;�4�9�d1���7�KF�� �������〯c9��)0�n�҂��vD��`�AuQ��/iNhz�-���H��<I��#���>Sx��U}Fx��NK�k����L�$N��8dM��}��F�J��7����:��_��n1w��:ٍ�;<PTң]�-e����� �7�H_�$N"�A��v���a��rnݞ������ŀ�
�MA�n�lx�[� �51RYw܆?��VT��!'MoK�&�9�:&B��)��*�X��*�.Oj�8I�Gƍ���gf�<o#�ޠ�����^��)����q��1���>����Ń�����:�&g�	W����O�v���b��4-���Tˠp���V�jy�Ru���s˴Χ��',l[k���p��
�ʔtb��bcZ����9Y�
+�s|`�1���>��"��m<t�11J"*8 υ@	�>$ًW�ENŃ�6oH���g�Ә���8�]?_*mG��WjIIo�<�.F����P�h�U�B�x2���ɣ2|�?����
�#2�+����;ng�3�Y*�Qg�P��MJ��cR���@�M.H+�ز�L苫ݕ����2�W�1}�D�m���{�F�
e����?-�G����w! ������ᩯIq�@J��`����	��eo���._|��Fװ~�r�)'iA���U�{�)\��9�p�l���̺��B�|�1����Lߨm�{i�H7�ЪQ���.��M;'�'�Ç%)���ԧ̄'V��M���a�d�ý!Bc�L�z+
�$uL_�`�~/�_�g(�Y[�fl'j�&7�#����@�C��,V*���eD������.̪��~ij�[���	�$��=d
�B�ȕ�I��"i�Ni���#R�>]|�OJ��_o{�I]���������L��ahI�3c�u9Q/6rj�V�YWCǁ��72ӗq<b}oή��Z��%�g��$�i��qI���xt��V��M/�76Ǖ ��/�>�-��RY�<y6����e	ԫ��+�b��������L��fGs�߱�n��|8
s�2;YF��?��N�Nn�c��%^���M��_2�
�G�*N9���4����/����ـ���C����R��$)Ո#�a2k{R�]�|SZ|��M��<��yE�&7�:[+�B/~��p>�|b���LEWU(�à���mdR�ȶr�ω�[s���>�Ne��)0�֏���.�Z����HxM( j8+�᰿Y��;���R��K;<+bE�M�7A��@�_j�������O�{J��?-�?��"�Da!�J�	i)m9q��'����|���Sj�����_�wT̋��n��@�T���;�HmF4��k�j��Kf�y �6�҈�����O����YKRX��:�?���\9oK�;��0|�"2ZvvM`͝�#&�P��*��~��p@ɖ����D�x���9D���2��n��'�a�,�#�r����l� �|y`��?D�<U� ��UU8=�����q�ܥq�$L��R�p�m*v��r��������'�)�OS�P*l�r��f�����)�v
p��̢*ڌ���]"��M�� ��#�<V���?o��9?K�'� ��(0�4j�Kb���NYb}�/�i2��HՊ+���ߏ��\����O��s��t� ,�C��!�VFN.G�l�4@0VJҪ�~Z�T?���oU�w�}p
&�v U�1�q�cF�W����f�H�䝓s�^ӿ�Z)	�Y��v�Ɛ� ��2�Z��Jp?�i�:�oC���J��X� "y)�<��DX��x����߰s�l.��w*�H
�I�� �����S�c�*@3)-�H`���_��rL�R�3X��b������lv�i�Z�M�5�X!Љ�-��1��v��5���cւ�����x,�x��'Rxm��f*l�˖2�1�)��i+]O�Gqhä�Vʂ�ΆY.W� ���r�l�	Pv�P�mr�`v���2f<Ɗ���/�h��O�bG���y�!P���&�5e��
-f��*#�E�u�pbM��!���C����;��˓g|E&W��g?+�>!������]"����	Z�B�^$�ɞ�:����*��@}ѓ��)�k"G�7����t���U�B�8�z@_��b2�ę���Hrj�En\���k����_K���G~��Z��T~\e�v��5k8!�����k��?�QF+52-���h�#j��o�~��W�8�������F�%y�dnאK�l��16}X���7h�##ݍ'�w�%��Eg�_a��eWZ�m<�P?�E�F�� �b�۩7��L<�t`��9q�E�:&��b�~���d�5��f\�Qm�9���GV	�;��sU�ch����Ǘ��?W�QmO`��� ��9�Y)����c�7�`��{5�l�D!��\RAs�<�M�~p4�ohQ��x �%��V5��l�4Fx��i�ŀ������lՅl�<7=h�Y2eѰFpxţm&��֪9���LǪ��E������E�;Gd��aHb	�y�����V�����I��= �͗2�Z���b�uT��٬Q=켸��;8P���[��\i�� u��-��(l��Vª���S:U��>I_N�V��'\�$g6Vg�S�1�~�1��æ�G�h�*��C���7í��������E�V�<���F])�B�ȝ���S$��RFKn��L�_VmdT�骆��^ �IΒ����� v�6[� C�ڦ�h����;���)VX�@�<�a�P��e̞Q5�)��nF~'Z�di���%f���4�z���{J�� h�=��S#;�ta��x����QH��ѧlW���3�l�|Vz���"f��@̎�2��������
�j#
b�ֿ ��K@�x�a�A!M	�Ҿ����3��j���eaH�2u�р�l�[>U��ݔo9�h_�S��!j܆C[�w8�P�c[�( i ��e�K{��[ڦ��J��e�aRs;��X���y�6��T`�N�'r�R<�;%F��$s�7�z
����S�B<Nw-���0� �̖I�y�wx��!��&���{�"���уE!}X�ƨ�a]��~����Q����*zN�!�_q���pk����֋��y������Q����.�!Ӕ g���cz��0XXK�\���Wآ���"�C���*�Kv�)�1�Q�n���8����5��Ai�n���].oO��m-��q�M���S#�L�G<�{��l�3E�X�6
	�K�A���X#\�+�44����~,p�RGAnq�4}SzDu�=ظ4l_	��Era"������G՘Gu�\�A�����b��^����0���a��ǲd~JL1H�������v�L9����@{9bT�_�%vQB����,�zy/S-w�v���H�ʼ��@ �1JЫp��Ϻ_ƦƬ6��l�/i�Y\~2"I��2��C(�d-D�Wx���ݾm�o9(���4ʹІ?�Ly�0O�� �� ��PZ:P�X7���n�4�#�:�}�L�:�k7N�ʂ����&������
A�}i�1��"�b�+�OB(O�<j��E�<&��5}���ڴ�\��\hW�fboW�Y�yI����˖ĂVk�f'���!��51�zΓ=M�fv���&j�a�U3�qn�v��B�g%{+ 7��"�ߣ��T ����Z�O֗�Α��O�'�C@둮�,s���[��)o -v[��ϡ��&w�S%o3�#;�,
�^n��/��!⊥���CJz����J�q�)����I�ތ	'��g��o��9��x�4NB� ysӔ i��dop>.t��z;�Q��{|���x������n�Re;�q@��f�8�Qhb n0�?����Uj*��&�p��	VR;��#l(�WQ���,b�H���l�/��U�n�e��W�z宿��z�r�E9N+�:��:o�&3^��o��)��V���h�s*�)pV(�1�)`|_��DHFWKD�m�:�FD9�Y����F�����<��&{�}10�|��bp���v%e�p����Y�f�=>k��4�D㵪5���2�l�J%O	�"���}47.�[1BڼtCz���/��ԛ��a�TGj�0�, Kmŝ�mEù˧�����s���r��ۈ.Ƹ�h�*պe<�CN�I��-GU��_{ -���r�*�g�3D�u�|�E�P"y��}���dC�����6T�ϛ��<)a���1ǚ��#P:l�5T^wbg����d�lt2��g�&�������e	Crv��r��L���I��/����\��~�:�]Wݧzߪ�G�o2�_d�W�����4e�T�7#V��֛V��X=X�j���@ʬ�m�^Jbxx�Z/T0����{����E߀���?���Er��3��,3bCv���
��M��
O��f!������QUJ�6w"	�u�y/ٸ�i��+%��L�Rsn���׍��Gx�]�������{�懈ſw!w�Z��nc�px�ȍn���b)�ۤ=�U���i�����o&��#�c�;��d��2��_�P�#.��0����  �r�̚�=A)%��~�;�2
�D�F9d4	�Al@SHc7Q'Xqa�f�<��f���&����1y��:Xz]:���&71|��A�PS�ufu�J�#�����Ye����b�[1�k�|�;S%M��o�BjQ�Qv��ղ�A%�(����M=n��q����V&��z@�xE���
�dAl,�?��q�^��w���U�X�ȷ�ǃj�Ǘ�[�kY�b$����}:�?r�������e��.�������&�$�X��P[食�9�Q���H�냅B�wȊ
��3�#���pY��O���n���o��.z�E{#o�ę jSFSԧdToE{�Ý�s
�cj��<|h<��`RC:#vn"ȂO���?:Q"�5%�1� 
�ڨW�F��1��N5���5?��H��>����~�$!��*�z�.�Z00�v�tW�Y-=��ih[�l��K'-6ؿ�JH{��/,�Z��ѭ����d~��+��t尨�=�߮��2��D�~5���LQF��(D3�,2%���"0���i��u�l�zWB�dT�}��y��C��Z����24��g%���YY�H�v�������b��K�[^`G_ �Ŧ��SS�p\��#'�n��M��?�"��{v-��}=AE�����?�h�@�&!�eA�N��I�
�w���\����b1�,��d����Jx�5��I�>gR�TX#�)�T��� �-d���a���h�-���xX[;�܂�R
�����֦��?ӛx.4�cW����C`�r�H)�$x��H�}J� <��^Ț�m���%��:qCvpB�#F�L#Y����@�D�o|�Jc{W����@�;m����X��O"|�q� >���r�è$�/��,�^=��/w� ��:���Au�x�_���SҊy9`��0bS-�$Eb�?=7�&��|
��J���z����<a��g�4��$��v��ci�r����׽�(R��!�����̽T�2T,���F�}-c��_�<�Mz1T>:�JC�!q�P��V�XHd���l��YU��.�"��O��з������6&2�`��iAd�[V'Ă̲����h��cچ�-�U���joW�_��sR~�0J�e��-6��w����.-z��Y�^��&֯R�K�!�Ҝ��S�8�,��:��k��S�KJӉ�����uN�,��(�Mz�I\l[�b�DGl�2ތW��1*er���R#�q�(ˑ����&y�6�2�u$9�B��Z���T�`�ؾ���F=0g��v�;s�&_S�d�f����R�)�}ap[1���<��>�K1GcO�~� �=Է�|�Yi�GBnY�~�֞��zpDZ��*Rѝ/\l���`U�t������1�_gm��6j��n���%�3�p�Yb��K�U�z�������اc��O+�N"������An]�-K�;vL�T���$������=�q�!����d�O��/��7$i�ڬOg�\H8�o#1.��o*��v��굯�,�D�[�A���)n:���6)ߧ�u�(T��+0�~��6gCc�R��Aɭ���x6k����5S���4�H�~`u��M:�1(��\�'T�JwRN5-�o� &�:�	��������ۻ�@>\���ݤ����EWy�i!����ώx12��,�tv��y��Qp�(�#n�1I�����#�������CnM��s�v��RYItuA5U�%Gd`�A��6<ϭ��A�����^���T�^�Q�ک����
�R��[l�r���b:�,�Mΰg$���kv6�� �Nr�����L�=�� O�����9�m�N���π3���nʈ*�l�ӈ��%�;A@�Ek���+� ��@^�Q7"y��H��i�f�>ߢﯥ�;��O�bB?��j��"��]�k����C�K����D��0	3�4��
��2	��d
I#z��t�����n�n�H4�J�'w��0ݳ�s�YjDFm*��z��m�n,<1(�bp/ރ7�A�?c���S9�_W V��x��g�=�ѷR���d;;ڧ�`�ٳ<qdq�;�8�Y�<��V��eZB	�mq�2@`K4+Z�i�ݯ�N�3'��1�T/r��ʼ�be_��TOz��F��W����� %$�)�;�=�8^^����$�l�
�_D�?��X�.�cVP��&�$���FPgS��wI������� .�E�T0����*����1A�F&��Ks�O��܋A��ߴ2~V�?A������ƃl����+ǌ^�����uG0��P$`_�>���߶���ݶ���-��wO���~@�P�"Ƞl�j��j�!�I�ߊ`,w�,>��� 7
��B,�O�VJ�����!Ds٧AO��������K�IJ͡��o�8ͷޖ�(e�������e�i�3�kߵeK���4+{g���UQ�$�p��� ΣG)y�';�8.��x���+� /�P�λ7�)�?���<[�
�3ү!LV�q�6w9np|�ߝ�g�qY��j�9~r�'��y�}�>7�&�H�؍1�K��D�
�! �9ᴑ��W9�]*-�����ĵ���Y�"6�1��J�gr\�r��-EŔ�f�p�K�5ù���AHl1��+0s �(G�ϯ��x������~I�iH
 /��	�=� � �5z���z��n��x�J[N�(�g5�'�\ �,�>w��<�V����OȬ�vQ�N��|HJF� }>��1�z�I�O�{�2jA�[ }�w�ܺ|C=��SAʽu|��2�-���:sy���¢[��q@R;��I�
|�VM|�c`�u�q�_{��з�!L"�X�c���t�8��m�=�� ����m"��sFVICC�������%� 4Qd��`��p�kk�'�J)n7Ÿ^�A.6��)Q�z���_ė.c%���`�m%gh/��Y;Z���3�����1���|Z��Gw��@o䖜4��`&�K���!�n���,�ٳ�Qa`����*��Q��z�a,\lUz���v�S!�A�RSC���&���B�y�3�p��O�^�~DJ�%L��[+�]�9�a��';�d��e4�)V:GE��+���DčJ�YG!�3g�m�1��(���l=�~Y���廦�o��=k8��9̇1�{l`}������m�^ڟ� |
WH]sv��h�=TNU���?�D\*�;o7-"!�\�� $�p�.�������y����(�^�4L�sl��>���dTR���	�wQD�[N��@Ϟl��'2���ׯ����p?��>��)�_��0�"p��B@���˼[ԁm�J�����v�?��p<�����s��z��5��*�}y:4���p_l0'�+(y	��M ��3m2��ei��w~g٭��e�.��]iK+7��'#n�"�|��ž�PiXrpR1�лD���R\G���S���V^��M�ޥt-��v�8�K��$@&��I�j�Y��r�9��&�L�GTy3l�V[ �z�L�p�Bǲ$.�h# Yo΄F�5���r�<���(������u2����3ޏ�[�q��_��
C��A'���͙e�ryq��(|�����l�[��m���JV��U@%X�a�L��察iyd�[��y����ܬ2F�w'��[������܁j\�W���3�5v�E�IC�s#��9s�M�z��,7*E��#s�#�Y$�M+P(6�@��竹�[W���%��O,��N���� � �P'�N@W˷��8N�	��n^k�e>�(6�΁(PMS��5/���b��4G\iFOٖ��3�)�KC��<3֎9?��H��=�iN��1W<�x���FK�/c�uSCE�'u�7U�Vz.Q )X�����ݝ��p�0�S�<�.k7�p@m����08�)��2)>�V�p|c�F�:ŋ}B�(�"�"�[����l]_�*���8��>gl��e�lQ*�sX!~��Z�8�Z{d�g&>x�qX1�g����#�����}�R�X
z��h[��� ,�$W}:���-I�0���Ul����n��0�%���F�hq)�2��
�˘w�W��&i��Dz	`}"~x)ኢ���Ӑ$C�*_�9k{&�N�R!a[t��)��� �VR����{f�
![���ar]Rͽ�aV�W���G���,>��!�q*� �$�����4��Z0�yE��ka��~	H&~�oг]�+�kﮢ�_����$��R��P��&�J���Z��ayʵ8����������j�T=�j�Z�Fw�^�q�nw�����D8�����>l�p0��%��Ύ��gD�r�w�_�]^e)��b����/ '��a���K��AKq�#�O��8N��1�o��ğy�b�V�I�L��YR�ã�b����~o�ٞ�p?L�*&2\�x�:�h��up�u���J�:�� �i2�w̅���	�AS
G��G����3p��q�')�E�I�I��6�R<��u�(���wO��H�xҠM�Z9����xkG�	6��8�ǌ=����{n��@q�@��27�h1�4D��\�R��%�3dm8�q:�V��m�gV�����U�SpT�l��b��&���X%�*&���8��7�[�N̡8�o�H��Y�<BGǮ7���o��k]8�9����B�h��,�xz:�;�I���p�@����LHo�f�����ie��}��!д�����H�BY��#��͖r�%�$�N}�X�  f��s@��ȴW�`�:��cjO&#���%��>Y�K���n��!�~��Jۖb<l�9��3^�����K�os�b$�|�swZ��O
8e�e-%��v�cx5�/E�4ᦛ��������#�2���4u�����./�oO	č���K{�EJ�lza]��N1~|����%zT�B�h���b���a�d�}�����}"��UMK�c���.}�#<|c����5
���eG5��$�A<$�h,����f�4��,Gf�7W����O�0h�����38͗��#�_��(kb>4��9$�+����)�=i+�Mݸ�eT�\�.�Vb�{%6<�v�*L�_c��ֱb���U[��1��n��ld&�X\�}�6
"�?�ӭ�V�:Q��\�O!�nC�a�E�"tܥ���=�r��p
�%X�t����Z��Rq�ݣ�+H�c����@G�Y=A �˖���������8Q��GL����W���c��gO%)�J��I͍_	�A�^�)��9m�J)�ΏPZ+�_���/>~h��Z�2u0ԡp�����&m����g�[�\�b�qtW`�&�f����uLP}��	��r�SY�G_�d�N���79���9�]���a�"\�s8[��i'K�ƾ���S7A��I$�g,.(�B;l3���_(�
�O�p�N.S��&�k��f�:�]W(��t��A7���&������@�wj���J���#�'���Mq ���D7���G�S����MU���S��"E

��=f��u.�Y�E��=�e�����"��f�;��k��!PB$9uV͖/��� ��R�����1փ��Ig�l=��M\ޞ�b��e��k�#���7�:ZvT�!{%�t�|��@��g3=�q����M�v��V�U�S�08���f6��j����3d�2G�,�/VJ�e�V�f9�s����'���~;^d��f�pUP;�H�+�z��m0mR�*l���P������z���-�����NLT��K��j��T��v6���8��] �c-g	(`B��K[P<y��7`v��ց��'�pM��ʏ~�M<"���2����\���3�)��e�(+�s��Q��GV̎����e�
.� ��Y��T�S�q����	�&���?u���K����N��ְa
`B1᫢�?HK�H��&{g��	Nr��xX[�N2x��������,����9�c�Kǻ�6�5�ǣ�M�*�;�;^�`/�3�Кx#��aY�� F�,h+�,�� �h~�a��o�<:+�W��&��p9LX������$�3�1t��F
��Nb��q.�؃�4� ���[(Y�6��Օk�$ŜbUqe���޿+q�9ץ�_��&��w�nה��1�A���M�6ґ���M_s�8:�`�U?���@]�!�L���8�;f�J��vGg0(d�?��\j�;���<�&�� �Ӆ+��|� }�U�$��=X��6Jr��|!��T���"�� �ӿwY���,.]'���;��w�����j��Do�ƅ��#������XK��;����@�i�^�7h�-V�8�,�bƋY��@������<f2�-I&]*{EZ�Ta0ЇE�=��-������7Q���]�m�`�וjŪ=�}�q4l1*XT2�<��O�[;����79l���!_$�MZEc�<��p�����R8F?H��aZ�L8��%a�D��n��݉g���ɒp��>��R���6E��_�c�좎�j.�J<̒v3j10'[�%����Jr��'����v�@���Ƹq�WS�;�2һ�Kg�ĳ�f6w�~�Y�ڰN�u�����dx\�(g�	Qը��#�ך����[����h��M��i���~;On�:�7������ߡ���>r$��S����#gg9�
}���5w6���1�Q+͍<z�R���bM�|���N��Cm-ظ_�4�R��`�cx��ȍ2_��:�ǹ(����Vzms[Yw���˔w��諷���
3Z��G�a�O ��^^;� FO����y�;<�sN��xe̽0�ej�ȵ�й�|�O���2�qy"�a�W��s?��A?#��3ġ*�(��fT�z�LeВW�(�R�	!\m���*>��4L�b��Vu:G�H���E=	`V��o�]ı��и?�����s�*�T�s��N ���(X.6�wI1b��5���V�����X���^���:��*ŗA=Ь A�Jg�Oj.29��L���vv�=�y������c�w�=sj�*���P���<6�.��}�yfV�c����l�����i�k���L�G��eY�Ɨ�M��̿���@�~d8�|0������h��x�p��r�0�>�VO�h8h6ujTH8�� ��M&ܼ�N���Md;I�[k�JF]���$_�=���*���b���Њ.!'�����y�A=�>�v�c�
�[��<H�9�P�Ok��u�I�{�辴J*>]\�8���}`���֮D� )i��e�̻'1��a�|�F�c�!��LM����M��sS�������Ү]�-��d�v�ܧ��,�|��"��
������B--[��UM���0��%�:uL2ݧ������lg&� (د:<(EJ|�)˪�ì��ST�K&���Fc�S��1HW}���^��n��E��t0$i<�Ǧ��;*�!k'NMs1"��MɃQҡ�71�p��s�׆��_"C� gA���^�+�I�<y�*�����.�w��F�e���/g���؋��н4U���,��$b��{w��>�_��S��%���ٙ�[Z`q��N��ͬ��ZJ�&k�'yâ@%H�M�D"�9�5�`����W�(O�F�E�x��c��L�t<�����rQ�+<��AM��j������d5��Đ���aŢeŬ��� q2:| mA��f�& |X���6N�2�影����@*�]���n���\�R�k�W�M�<&���jy!4N�'.�{�"����n�+!%��yݾ�V�n^8�4��\��&}���h�~N,	�:�K.���8rg��N���&y]Ƹ2-z���UT ���R��
zN��	yŞ^�ⲻ�6x����)9�i�I����l2�|d�W�'����<W߰�͒�b�R��HD�䖆K�l*$��i��H����z�F�xa�q�Z}��:�|���xʒwJ/��tH	�ʹH{e
,���т		���p���{.�W�J��}^����.JOv&��o6����Ɣ`IV�`�	fb8��TM��N
���Z��-�
�8��o���Ӛr��Y��fX-g]�b?�g02 P=X#Q���ъ"�#��s�39�G��		��N���DJ�pL�]|e�N�����\�nस���N��R5�#M��q�JWR��.���ڵ�#1�^�=lC���c�:�^D��Wo~��6�p����9��<_��|�xƚ*[kc�����$&�����	�
90���%Td\����4�l��s�8	e����(�M[Ǘ�ˠK�](�f��Qh����O�ZB$`�X.��4E#a���,J����o}�a��s�k�nTƖ�4���aO8+3Q�z��H��?�e'{T7��=#m/Ih뽢�xp�8� ڥ8�[yHB�#�r�������yI�;s��F����Y+�e��"��.�#ߑ�P>��c�ލr�)��b�0���z2qUwQۻC`}�ۀ%I\%$�w�V���1�C􍽰��L,�cw��R�5edm#�E2G�)��F�s���'*��pa�J\Pmt��OM�$3�� �M;� ���"��+�3�'�w���qK��������$_4���ݒ��)�r��X������WϷN8��3���Eѿ�a��t�7�f4(z~��S�͙������	ʝ�cG�g��!q��{AO�Sø�Y.�"ۿS�d�B�o��/�v����S����񚐭��MZjX$����n��C�j�Z��X�u�{��:1��Q�WY����U���/"q�����5�A�Ce��kb/���8��TM�H6�X�O��x�`�O�a�;LU�o��bq=.�����~uO¸���ǧt%R`&��j'b�&<- @j����S��32�0��j�¨iq����Pd�V�R��_����9
E _zB��X��(EQ�֛U�j���$Vcj����!y
���,�X�6�jFV2��g��&�7�'`5��`���oy�Y�*��|�Q
!�#"�:�s���n�%���1;�[5�@c�q��!`x�L��M@��'����[W\���LT��4r��T��f���vlSd{ݨ��Q1#��_� ��^qM~W��[�O19�aT-[N�m���yKn�Y>��@���#ؑ���k����m����Y8H��I���ВTm�8f���~@E�����R��\_�#�.j�66�Z��Ew��"�(П(+�q�]I
W�D�Ԧ$�>�����8���֙��_�Mь�ʤ�z�_ޯ���c�v�����{����CE����M~�/����'<Ņ~��;��,��)�����BT�VC��(�N�\�9� ;���5h�T�7�_�@pgm��7��$e��H�O|��B�3?L9bO mp�����	X�+%ź�Wxp��1�M��u�@��S��s6Z�Bh�-A;)$�]�� �a�GlU����ը��?X�bK��C5��p�Fs�L/��c"H$��}��u�}��2�My����]P0�}�2�m�T�~�	c�u���@��P�xBI^�t�j��q^��H�e�l`z5gPV˼�^Vuz�~���|��#G��� ����*������`ڴ�7���2�ErbC1�:Es����~�ks~�0�2��k�9ZJ~u��;E�~�rE� ��	�ǋ�I>�xQCLV�����KZ�����L�)7l#����_A��1�
4�		,��:�t1�8��\����M];el=�x5����S���k쒆?'i�+�f�_��>�E���3�����%��ޜ6��J�>j��H|b�ѓE�K�����Ӷխ�ϒ��1K��+�r��+&�a޳F�-�uQv�'3��[SM]mF��?a��rs�P�8A�9��"9��@pK ��W3�"�e�c���j�5��"B��:��q������=��%��?�uyZ��*m/�^�߮��w(g�#2�S>���\S�{�g���"�e���)�F�u.�TVu<h� �1˓a��vj�ZL�ȍ�e��d@`*'
���5M��{��SNyP�� ��K������0��Xb��B*]Rbc�0G	�'/N��o���0��X�õ@ 	%���"��)�I�*��,�����Ś��|hM��Y�ɛh45��b�n��@5�Ď���v���_aU���Qv1n���eD2�7�2sBR}����dA�E
#�P>�	D=E��Y&R'��Iiu/z�+PG0�-	h���b����Y��b��x]�����0��
Ka�{Cp�i���� g��߭�����5���D�}Z�R���l܊h��}y�㪌��7W�H�.Q�
V� ��g&s��'S���O�C�J��ysN�g=) ��Ž+�Rb�����Y����BU�6�:�:���A"�G�,�� ���N��h�>$�ff e�1�tr�$�Q[����m��S(69��j������Q�y�m�4$L�ܔP"�LM����C(W�<��P(ݷ�G�ry�+�"4>���~Y����y%��>(�����|�}�qSFr�㢩��3"�����d�,����k��6?6��`��+���Đ�,��n5���y�$��!v��ƜT\0<����A���(�tVEC�0����u^��K&-�-���t��~�)�����(/�{�t���:Ր�KW��Y6`�Ɨ\��i)�+������^��zl���t�b�Q��Q<���.��Q��{h��,LDU�$�X+�����=p�-)��d+Y��s�.���>��a0\���'�'������1��d�Ղ�W[A���ؒ�V3dyc�/��L[�Kn^] }�V�n����wD+Ӷn;)��+��yQR�%��s�)��g�����1��`�G>Ɛ���?����{�zQt	N�s��Z4�}�Wp�e��0eI��κ�c,���;g�W���)E`���`-�����w}�b���t(�1��Yu�vш�d�hGht ��GM��	��s$��LK7�i�w��~F��=���VL�?Э�`�z�
�n�D]w��5���Ȥ�H������Q��\�]�Q����] �w8L:�Q_�
d�D��ȉ
e ����_;�5�R�s�Vkr��*�&[�IJ���${@{���!4�c��_�og��M�֏^��te��d�+�eL�ɒ��梒%ݠϟ.%�UQU��t�6.���}z|-
��W��aW8�m{Y�j�u�w�Z�'ST����+s�0e�Х��^Ly�l���4���|�0�a7)a���O*j�9� �w�Z��=��d���7���>�j��Ƀ�뮟=Q+"��*]& �4Z�熕%Q��R�TQ��<�nR�ч/���,� �]8}s2f��{�������]̰/��"Yɷ�pL:�H3�F���w<F>=���k	vs3���qzg"8�A;2N�K�	�����Ņa��wܿ0�&q����T�^.Py�5���R%���\f}�d�9��ő�*�|�#�;
&懚��<W��~�겶
�%�3�ܴ�B���-M��eA���p�iy@#j��r�X�^��Y�԰�NN��)���6��+�BEu��T�0�&�Hh�4������nj�)�W-����V� I&��$���7お���%���lT��/���F��6(�n���_�sl}�����ߕx`$�N޹ԥU�o�J@�w�A����`�A��S&[eŦǟ���� �h�_�a�|t��3���a�
�z�i=�}%�N�Sծ��ս�$w�(�3s`/u^�P��.�}��~&�0��ނc׭�mi�(�u�c���<S`�"}�����W���I[e��u�o[��m���|. :�o1jdS���i��%�p� �.;��e�j�d0�^C%Fv�<ԩ��0j�"�#�2�a=�a���9�T�-��>���]��_.�M�G���Es_��?���%��2h�Jq�h�-:��F��|�W��ӿ�/�/%p�)��'!!��fȼytm�vTǊk��AZ�6D�>�~�
�ю��Wz��F��Wn��vz�ͷM�s�ui�1�ǻ)��7o�J"~���㠇Q�X�m ��[L!>j�/1����E��jSׇ��CИ��[!�8�*n.	�y5���N��׵9]�+�)�9k2�Rrn�ݕk��IS�=��`��zg����F��x/-j�G��f7�9m{����i(�$���!��Tc�lG��ǰ(�ө�в����|k�����#�*��~�u��I7�n�<�:�u3��V�(�U�x�N��K�KI�*�1uF�D�| ^/Q��������뺘Ͷ��}���s�=D�hT�R)���7l�\����B/�����Piv��i������ܱ]�+Y�v6��Q���u������>����G�A���
^b�.R�I������(���]mEb*���.�~���[!���+��dA�Lv0k��#���-ɹs���%�}�V����%s���u�u@��O����x<4��y��:�=-�s��_�$�v���&�O@nv��e����:6��CT�.0X�Ӈ�EʢH챸�#�mg-��q�H��l̊�ir2[�"�n �l2?�P|XVo7�k��Ŵ�a����������)v�FJ93R�li�+�mG�)��z��L�J(I,�
�����%x��M��-LhE��ŧd&a���a"�p�	���~�	�΍b�A�%��2��*��]��0�XD�g��@S}O��a�ܼ;6�6���UZ(ҧ>��9 �4��M!6'I��m��2���wI�k3�q��A��e����/�ξz���uT0_���"���\��^�ӘYK���s����t�d<��w���i��[��bvV�G5��71�k�\/+\l��kbR�x�p3���%kf��9)%�I�b.z��M�^��[��Ş%R�~��?s��+����D������EGE�r��AV�q=4���w��*���tm�u�$'��_�1jZ߶b8�u�9v��A瘱���J��>�`Ms�������R}�F�谓`��FN�_i���lVY�<���[��a������7&����ޗ���H�K����Ku3��PRK���_"9Q���
I��]y�,��!��x���������uD��ͅ7Q7��.����6c8)-d@����۳����y����$x�D_�#ή�O�Q����y<ݘe �� Jb��ج.�T_�*�U�]��/|�J6���i�*a�=�=�aFJ�.�*F`����i���"��+tW�����M*6u�{ڃV-�tA������k����{]���	��L}M"�܌�Lp�Uٶ�R�w�,�~�JIgK�?�R��a#q9O� ���2�J,eO#�3f΢�<�i�×B���g�p2xėd�9�v4�O�����g�h�3ɥ�O����x�C�4iϴ�{ ��!�7
	�Aܻ2��tJ���}� ��9/�y)��ĤJP�9�؊���:�J��T��};��-[oN���y74�]`M��2ze�MI�w�A��͵g�3�2�z��n��5�$�f�����(�Ԫ�>9,�'/~�BK8F�&�6ɲ�>��Зj �*��Q͝w1�O5��'߃ÛE� �i��ڣt��p�ۄ�Q��A�xV,#LN�w�s����1eX ԁ�R��^XԬwBJ���v��5i�z��}���M����~��̵�7`��4\�4ݬ���M�Iп):�W��2���s@�Y�j����R��������og4�����j_]4�*]�n���w�d�qB�4�&���hLi�\'TB�����=�J��;�=i�Q-�(1;'�ܴ��Bf��y�$a�&�G�������j�R"�F7�h�~���j��3o�{ou��J�J�F3C�RB��ZQ"�.^EY���fC��ؽ�s�S���v�
o-�Y�&���H��٘z��Z|R3U.M��8_�4�!X-1&dEd:�)�ef�Dr��|�v�]�k�|�8���Ȓ��& |"8�DIs]���}~g�kY�zo&� [9�ǖ�E��A�8Ǘ�r6�27�k�y�a
	uKM�s�ް��m�FޯR,> �v�q�^V�@�9�) k�ׁ�����W͛����9d�|a����_w�F���yR�|]���G�_��(�.^	Il���f�S �����o��S]?�HJQ�<�
 4i�Q�B��?�\.0j~D�m��H.��h˝si�4I�(�%��X���d�}��� ��F��	�H��+�
cy��1��x���WqR�Τ'�#�,(�'�1���$�f��#�v�-�l�����&�G	f���logr�{B�q�3rZ���d��>,=��2�\oa�tm�=�3�\���x����s7�t����Gmn��(3��3j3�K�5��2mTݨ@��1E�-�Q3�����X"����a�i0�S&���C��K�/���n�`R�V�"��m�|�U9���{8Z���������y������roR���Aƌ���҆yM��:Q�J`��`ICۗ�+�&%�XMĜ��Y&��M��f �b�S����t���e3U�5�͝�r,"P�4�CP��L�����y��E�(��J?|�gvJ�SR�$y.oJQa���{NNs�*�a͕��f�f�}�+4�뇦�5h;dIb\�-�T���V~� ��e�:�_y�g� :��di��=�%�&������'Ȫ�8�k@RC��8���U�������&y`�F��^���3+!��C�ΰ��4r]fK��^��'6݊� �6БP ��4K�3�����
�<HXD6e������2�N	���5�|$�" @��q�zqG�ru����U� ���L�o����7x
 p��sI�&���XtȪ������
�i�Ś��8�/�(E��,a�Ӽ�lJxK��T43w�ϙܵ�����y�hpׇ�@�އ�=��i�-1��t�O���N�k�5gp��g��S��<����i��D��N�w�K�b�Ύ&0����Ab�~�*�Yo���2R��1;��]���A�hlZ5.IM�7�H�Q�Jаq��,����7T�m�O!�lGb\��*�K(��'�뢱����$�@Q�گ�əNDgx���ܯ2��ec�k��κW�X)��Ǩ���o��<ѱ�ޣ�$쪰����3S��͚z�����u�p��DK��hR�r�q�	��G�_{�\|.Iu�=J�۾�`O�]��O��-䎢�C]�v�}N�J(�N�~ꚴ�l.eh�7� `��U�VBvf��Z�j=W�u����xMpLMس��FN���G��t[�c�RW�z��\�?vQ�R p�c^�?նm���b���Il�j�j_�i?�������g7���B�Ư�(�!љ�(L�=+��4Do �T6l5ӯ�����D�&��jt�&��tz���}?hD�a?O���WyG�(`W
�[��'�6�y9��_�S��͠&Xt�:�)(�p������<�nx�[�C>4����v�ت�>���� �������B�[�(�BH�}�ȩ��V�A��b��� 4Q���s	��r��	.�Ȑ2W>���)<f�2�  �K$H�?�T�i�~�/�3���5����j��v�l�����e,R��I����n��^?)�V�����	�>}��E��5�iU�<�<���q$�J�+�7�op�{����Y
��qL/'�W�vi���	3��y�!^����o�	R�e瀿�j2����A���u+�Ig��>�D[K�"�=9q��a�|�K{�*\�sH��ҋ�n|�4;�>4NjE�!_��D�O��i���e�ϥ�d�"ޝ!7~fUA��E��
A/L�����L�b%o��O�ͷ����^]-��Ø`���JC	Ǌ��!�b��
'�̅t��X�Î-e��e��5���}�ތ�1��71g�=���[�?�Ϭ��Ij�Lh}�Й�J\q�jOՂ.B��c�^�P�*���R0��D�y �^3=�[������%���r��o��[� �8˺K�T�*C�a���\a�4���*y>:��Y�">Q��6�e�!���HM-t�b��E�~Ha0x׈>�f������K5+�zN�:b�`"=5���X�k[cW�!Z���<z�󸘀�Ɛ�:6:CO&�ט�4N�#K+�Z�{z^�H=��h��S�tq4L�*ʌ�otk�!�:LM۩	M�<sg�qO�Ω�B�~wd�/|�yuVn�aK��;zg�B�1�xТ���k!��}�i[� Y*
�W����f�H�qf  �P�-=�@�(�7����4bʶ7�G�����"k�I0̴>���h���FD��l�cC<1�/`������L��b�Ս�B���IQ�-�\�c�(;�q��I����ƍ4U�z��B{�#>C�md��H�sG)�N�����7�T������2$���S�A��冝�o�:w9�K��Z��i�"Sh ƜP���nY�nx�O�>��h*�;ׅ�mݱ%�т�@:
�[�h����rw�]��珹�*�����P���Ϲ��J� y\J�Z�����iY�J%��T����'IY�C�xfһ^I+9�n!�@��� fvk��_
xV��iF����#��=�ҩj&Q>��M��>��Ezc,.]��-X��Qg�?���KC�q$>��O�=���Q}<p��TM�}c�3�,�]����#4�O���`ٸ�q��rǔ)l�r�{��:ܪp2�X�?��!�>Wj�������M�o�"&��f�����ϙu�gU��Ս�S�+_��;`��D�8�'�����DA��5�WQ����6	�l���3�R�3|̷:D�zj�:)�nk���n�;(?(Lo�o����WM!���dO ���� ^:�Vx�=�rp�*��ml��Rw^�O��J�~=��\$<[ɚ��#҉޸Ź)��u�K�u��Z���R��	Z*/jrZ������@mb����(nʍ~����lSK�����<9"�¬��)���j���t;k���VS����{��<ҮW���@9�u{�f���m[)������s*��[9
��T3E��O�[��&F������Э�H�y)���!#�e�L�cv�u��l��f�j�$#�GR/>�ώ�|F1�q�6��l�ȏe�$