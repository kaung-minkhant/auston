// DECA_QSYS.v

// Generated using ACDS version 15.0 130

`timescale 1 ps / 1 ps
module DECA_QSYS (
		inout  wire       audio_i2c_export_scl_pad_io,              //                  audio_i2c_export.scl_pad_io
		inout  wire       audio_i2c_export_sda_pad_io,              //                                  .sda_pad_io
		output wire       audio_reset_n_external_connection_export, // audio_reset_n_external_connection.export
		input  wire       clk_clk,                                  //                               clk.clk
		input  wire [1:0] pio_key_external_connection_export,       //       pio_key_external_connection.export
		output wire [7:0] pio_led_external_connection_export,       //       pio_led_external_connection.export
		input  wire [1:0] pio_sw_external_connection_export,        //        pio_sw_external_connection.export
		output wire       pll_audio_clk,                            //                         pll_audio.clk
		input  wire       reset_reset_n                             //                             reset.reset_n
	);

	wire         pll_c0_clk;                                                  // pll:c0 -> [irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, jtag_uart:clk, mm_clock_crossing_bridge:s0_clk, mm_interconnect_0:pll_c0_clk, mm_interconnect_1:pll_c0_clk, nios2_gen2:clk, onchip_memory2:clk, rst_controller_002:clk, rst_controller_003:clk, sysid_qsys:clock, timer:clk]
	wire         pll_c1_clk;                                                  // pll:c1 -> [audio_reset_n:clk, irq_synchronizer_001:receiver_clk, irq_synchronizer_002:receiver_clk, key:clk, led:clk, mm_clock_crossing_bridge:m0_clk, mm_interconnect_1:pll_c1_clk, rst_controller_001:clk, sw:clk]
	wire  [31:0] nios2_gen2_data_master_readdata;                             // mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	wire         nios2_gen2_data_master_waitrequest;                          // mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	wire         nios2_gen2_data_master_debugaccess;                          // nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
	wire  [24:0] nios2_gen2_data_master_address;                              // nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
	wire   [3:0] nios2_gen2_data_master_byteenable;                           // nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
	wire         nios2_gen2_data_master_read;                                 // nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
	wire         nios2_gen2_data_master_readdatavalid;                        // mm_interconnect_0:nios2_gen2_data_master_readdatavalid -> nios2_gen2:d_readdatavalid
	wire         nios2_gen2_data_master_write;                                // nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
	wire  [31:0] nios2_gen2_data_master_writedata;                            // nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
	wire  [31:0] nios2_gen2_instruction_master_readdata;                      // mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	wire         nios2_gen2_instruction_master_waitrequest;                   // mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	wire  [24:0] nios2_gen2_instruction_master_address;                       // nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
	wire         nios2_gen2_instruction_master_read;                          // nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
	wire         nios2_gen2_instruction_master_readdatavalid;                 // mm_interconnect_0:nios2_gen2_instruction_master_readdatavalid -> nios2_gen2:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;      // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;   // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_audio_i2c_avalon_slave_0_chipselect;       // mm_interconnect_0:Audio_i2c_avalon_slave_0_chipselect -> Audio_i2c:wb_stb_i
	wire   [7:0] mm_interconnect_0_audio_i2c_avalon_slave_0_readdata;         // Audio_i2c:wb_dat_o -> mm_interconnect_0:Audio_i2c_avalon_slave_0_readdata
	wire         mm_interconnect_0_audio_i2c_avalon_slave_0_waitrequest;      // Audio_i2c:wb_ack_o -> mm_interconnect_0:Audio_i2c_avalon_slave_0_waitrequest
	wire   [2:0] mm_interconnect_0_audio_i2c_avalon_slave_0_address;          // mm_interconnect_0:Audio_i2c_avalon_slave_0_address -> Audio_i2c:wb_adr_i
	wire         mm_interconnect_0_audio_i2c_avalon_slave_0_write;            // mm_interconnect_0:Audio_i2c_avalon_slave_0_write -> Audio_i2c:wb_we_i
	wire   [7:0] mm_interconnect_0_audio_i2c_avalon_slave_0_writedata;        // mm_interconnect_0:Audio_i2c_avalon_slave_0_writedata -> Audio_i2c:wb_dat_i
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata;       // nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest;    // nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess;    // mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_address;        // mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_read;           // mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable;     // mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_write;          // mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata;      // mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                    // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                     // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_read;                        // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire         mm_interconnect_0_pll_pll_slave_write;                       // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                   // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire  [31:0] mm_interconnect_0_pll_audio_pll_slave_readdata;              // pll_audio:readdata -> mm_interconnect_0:pll_audio_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_pll_audio_pll_slave_address;               // mm_interconnect_0:pll_audio_pll_slave_address -> pll_audio:address
	wire         mm_interconnect_0_pll_audio_pll_slave_read;                  // mm_interconnect_0:pll_audio_pll_slave_read -> pll_audio:read
	wire         mm_interconnect_0_pll_audio_pll_slave_write;                 // mm_interconnect_0:pll_audio_pll_slave_write -> pll_audio:write
	wire  [31:0] mm_interconnect_0_pll_audio_pll_slave_writedata;             // mm_interconnect_0:pll_audio_pll_slave_writedata -> pll_audio:writedata
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata;      // mm_clock_crossing_bridge:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_s0_readdata
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest;   // mm_clock_crossing_bridge:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_s0_waitrequest
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess;   // mm_interconnect_0:mm_clock_crossing_bridge_s0_debugaccess -> mm_clock_crossing_bridge:s0_debugaccess
	wire   [9:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_address;       // mm_interconnect_0:mm_clock_crossing_bridge_s0_address -> mm_clock_crossing_bridge:s0_address
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_read;          // mm_interconnect_0:mm_clock_crossing_bridge_s0_read -> mm_clock_crossing_bridge:s0_read
	wire   [3:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable;    // mm_interconnect_0:mm_clock_crossing_bridge_s0_byteenable -> mm_clock_crossing_bridge:s0_byteenable
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid; // mm_clock_crossing_bridge:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_s0_readdatavalid
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_write;         // mm_interconnect_0:mm_clock_crossing_bridge_s0_write -> mm_clock_crossing_bridge:s0_write
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata;     // mm_interconnect_0:mm_clock_crossing_bridge_s0_writedata -> mm_clock_crossing_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount;    // mm_interconnect_0:mm_clock_crossing_bridge_s0_burstcount -> mm_clock_crossing_bridge:s0_burstcount
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;              // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;                // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_s1_address;                 // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;              // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                   // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;               // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                   // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_clock_crossing_bridge_m0_waitrequest;                     // mm_interconnect_1:mm_clock_crossing_bridge_m0_waitrequest -> mm_clock_crossing_bridge:m0_waitrequest
	wire  [31:0] mm_clock_crossing_bridge_m0_readdata;                        // mm_interconnect_1:mm_clock_crossing_bridge_m0_readdata -> mm_clock_crossing_bridge:m0_readdata
	wire         mm_clock_crossing_bridge_m0_debugaccess;                     // mm_clock_crossing_bridge:m0_debugaccess -> mm_interconnect_1:mm_clock_crossing_bridge_m0_debugaccess
	wire   [9:0] mm_clock_crossing_bridge_m0_address;                         // mm_clock_crossing_bridge:m0_address -> mm_interconnect_1:mm_clock_crossing_bridge_m0_address
	wire         mm_clock_crossing_bridge_m0_read;                            // mm_clock_crossing_bridge:m0_read -> mm_interconnect_1:mm_clock_crossing_bridge_m0_read
	wire   [3:0] mm_clock_crossing_bridge_m0_byteenable;                      // mm_clock_crossing_bridge:m0_byteenable -> mm_interconnect_1:mm_clock_crossing_bridge_m0_byteenable
	wire         mm_clock_crossing_bridge_m0_readdatavalid;                   // mm_interconnect_1:mm_clock_crossing_bridge_m0_readdatavalid -> mm_clock_crossing_bridge:m0_readdatavalid
	wire  [31:0] mm_clock_crossing_bridge_m0_writedata;                       // mm_clock_crossing_bridge:m0_writedata -> mm_interconnect_1:mm_clock_crossing_bridge_m0_writedata
	wire         mm_clock_crossing_bridge_m0_write;                           // mm_clock_crossing_bridge:m0_write -> mm_interconnect_1:mm_clock_crossing_bridge_m0_write
	wire   [0:0] mm_clock_crossing_bridge_m0_burstcount;                      // mm_clock_crossing_bridge:m0_burstcount -> mm_interconnect_1:mm_clock_crossing_bridge_m0_burstcount
	wire  [31:0] mm_interconnect_1_sysid_qsys_control_slave_readdata;         // sysid_qsys:readdata -> mm_interconnect_1:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_qsys_control_slave_address;          // mm_interconnect_1:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire         mm_interconnect_1_timer_s1_chipselect;                       // mm_interconnect_1:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_1_timer_s1_readdata;                         // timer:readdata -> mm_interconnect_1:timer_s1_readdata
	wire   [2:0] mm_interconnect_1_timer_s1_address;                          // mm_interconnect_1:timer_s1_address -> timer:address
	wire         mm_interconnect_1_timer_s1_write;                            // mm_interconnect_1:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_1_timer_s1_writedata;                        // mm_interconnect_1:timer_s1_writedata -> timer:writedata
	wire         mm_interconnect_1_led_s1_chipselect;                         // mm_interconnect_1:led_s1_chipselect -> led:chipselect
	wire  [31:0] mm_interconnect_1_led_s1_readdata;                           // led:readdata -> mm_interconnect_1:led_s1_readdata
	wire   [1:0] mm_interconnect_1_led_s1_address;                            // mm_interconnect_1:led_s1_address -> led:address
	wire         mm_interconnect_1_led_s1_write;                              // mm_interconnect_1:led_s1_write -> led:write_n
	wire  [31:0] mm_interconnect_1_led_s1_writedata;                          // mm_interconnect_1:led_s1_writedata -> led:writedata
	wire         mm_interconnect_1_key_s1_chipselect;                         // mm_interconnect_1:key_s1_chipselect -> key:chipselect
	wire  [31:0] mm_interconnect_1_key_s1_readdata;                           // key:readdata -> mm_interconnect_1:key_s1_readdata
	wire   [1:0] mm_interconnect_1_key_s1_address;                            // mm_interconnect_1:key_s1_address -> key:address
	wire         mm_interconnect_1_key_s1_write;                              // mm_interconnect_1:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_1_key_s1_writedata;                          // mm_interconnect_1:key_s1_writedata -> key:writedata
	wire         mm_interconnect_1_sw_s1_chipselect;                          // mm_interconnect_1:sw_s1_chipselect -> sw:chipselect
	wire  [31:0] mm_interconnect_1_sw_s1_readdata;                            // sw:readdata -> mm_interconnect_1:sw_s1_readdata
	wire   [1:0] mm_interconnect_1_sw_s1_address;                             // mm_interconnect_1:sw_s1_address -> sw:address
	wire         mm_interconnect_1_sw_s1_write;                               // mm_interconnect_1:sw_s1_write -> sw:write_n
	wire  [31:0] mm_interconnect_1_sw_s1_writedata;                           // mm_interconnect_1:sw_s1_writedata -> sw:writedata
	wire         mm_interconnect_1_audio_reset_n_s1_chipselect;               // mm_interconnect_1:audio_reset_n_s1_chipselect -> audio_reset_n:chipselect
	wire  [31:0] mm_interconnect_1_audio_reset_n_s1_readdata;                 // audio_reset_n:readdata -> mm_interconnect_1:audio_reset_n_s1_readdata
	wire   [1:0] mm_interconnect_1_audio_reset_n_s1_address;                  // mm_interconnect_1:audio_reset_n_s1_address -> audio_reset_n:address
	wire         mm_interconnect_1_audio_reset_n_s1_write;                    // mm_interconnect_1:audio_reset_n_s1_write -> audio_reset_n:write_n
	wire  [31:0] mm_interconnect_1_audio_reset_n_s1_writedata;                // mm_interconnect_1:audio_reset_n_s1_writedata -> audio_reset_n:writedata
	wire         irq_mapper_receiver1_irq;                                    // timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver4_irq;                                    // jtag_uart:av_irq -> irq_mapper:receiver4_irq
	wire  [31:0] nios2_gen2_irq_irq;                                          // irq_mapper:sender_irq -> nios2_gen2:irq
	wire         irq_mapper_receiver0_irq;                                    // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                               // Audio_i2c:wb_inta_o -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver2_irq;                                    // irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                           // sw:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver3_irq;                                    // irq_synchronizer_002:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                           // key:irq -> irq_synchronizer_002:receiver_irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [Audio_i2c:wb_rst_i, irq_synchronizer:receiver_reset, mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset, pll_audio:reset]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [audio_reset_n:reset_n, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, key:reset_n, led:reset_n, mm_clock_crossing_bridge:m0_reset, mm_interconnect_1:mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset_reset, sw:reset_n]
	wire         rst_controller_002_reset_out_reset;                          // rst_controller_002:reset_out -> [jtag_uart:rst_n, mm_clock_crossing_bridge:s0_reset, mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, mm_interconnect_1:sysid_qsys_reset_reset_bridge_in_reset_reset, onchip_memory2:reset, rst_translator:in_reset, sysid_qsys:reset_n, timer:reset_n]
	wire         rst_controller_002_reset_out_reset_req;                      // rst_controller_002:reset_req -> [onchip_memory2:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_003_reset_out_reset;                          // rst_controller_003:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, mm_interconnect_0:nios2_gen2_reset_reset_bridge_in_reset_reset, nios2_gen2:reset_n, rst_translator_001:in_reset]
	wire         rst_controller_003_reset_out_reset_req;                      // rst_controller_003:reset_req -> [nios2_gen2:reset_req, rst_translator_001:reset_req_in]
	wire         nios2_gen2_debug_reset_request_reset;                        // nios2_gen2:debug_reset_request -> rst_controller_003:reset_in1

	i2c_opencores audio_i2c (
		.wb_clk_i   (clk_clk),                                                //            clock.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                         //      clock_reset.reset
		.scl_pad_io (audio_i2c_export_scl_pad_io),                            //           export.export
		.sda_pad_io (audio_i2c_export_sda_pad_io),                            //                 .export
		.wb_adr_i   (mm_interconnect_0_audio_i2c_avalon_slave_0_address),     //   avalon_slave_0.address
		.wb_dat_i   (mm_interconnect_0_audio_i2c_avalon_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (mm_interconnect_0_audio_i2c_avalon_slave_0_readdata),    //                 .readdata
		.wb_we_i    (mm_interconnect_0_audio_i2c_avalon_slave_0_write),       //                 .write
		.wb_stb_i   (mm_interconnect_0_audio_i2c_avalon_slave_0_chipselect),  //                 .chipselect
		.wb_ack_o   (mm_interconnect_0_audio_i2c_avalon_slave_0_waitrequest), //                 .waitrequest_n
		.wb_inta_o  (irq_synchronizer_receiver_irq)                           // interrupt_sender.irq
	);

	DECA_QSYS_audio_reset_n audio_reset_n (
		.clk        (pll_c1_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_1_audio_reset_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_audio_reset_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_audio_reset_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_audio_reset_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_audio_reset_n_s1_readdata),   //                    .readdata
		.out_port   (audio_reset_n_external_connection_export)       // external_connection.export
	);

	DECA_QSYS_jtag_uart jtag_uart (
		.clk            (pll_c0_clk),                                                //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver4_irq)                                   //               irq.irq
	);

	DECA_QSYS_key key (
		.clk        (pll_c1_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_key_s1_readdata),   //                    .readdata
		.in_port    (pio_key_external_connection_export),  // external_connection.export
		.irq        (irq_synchronizer_002_receiver_irq)    //                 irq.irq
	);

	DECA_QSYS_led led (
		.clk        (pll_c1_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_s1_readdata),   //                    .readdata
		.out_port   (pio_led_external_connection_export)   // external_connection.export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge (
		.m0_clk           (pll_c1_clk),                                                  //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                          // m0_reset.reset
		.s0_clk           (pll_c0_clk),                                                  //   s0_clk.clk
		.s0_reset         (rst_controller_002_reset_out_reset),                          // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_m0_writedata),                       //         .writedata
		.m0_address       (mm_clock_crossing_bridge_m0_address),                         //         .address
		.m0_write         (mm_clock_crossing_bridge_m0_write),                           //         .write
		.m0_read          (mm_clock_crossing_bridge_m0_read),                            //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_m0_debugaccess)                      //         .debugaccess
	);

	DECA_QSYS_nios2_gen2 nios2_gen2 (
		.clk                                 (pll_c0_clk),                                               //                       clk.clk
		.reset_n                             (~rst_controller_003_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_003_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_gen2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	DECA_QSYS_onchip_memory2 onchip_memory2 (
		.clk        (pll_c0_clk),                                     //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req)          //       .reset_req
	);

	DECA_QSYS_pll pll (
		.clk       (clk_clk),                                   //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),            // inclk_interface_reset.reset
		.read      (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0        (pll_c0_clk),                                //                    c0.clk
		.c1        (pll_c1_clk),                                //                    c1.clk
		.areset    (),                                          //        areset_conduit.export
		.locked    (),                                          //        locked_conduit.export
		.phasedone ()                                           //     phasedone_conduit.export
	);

	DECA_QSYS_pll_audio pll_audio (
		.clk       (clk_clk),                                         //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),                  // inclk_interface_reset.reset
		.read      (mm_interconnect_0_pll_audio_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_pll_audio_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_pll_audio_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_pll_audio_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_pll_audio_pll_slave_writedata), //                      .writedata
		.c0        (pll_audio_clk),                                   //                    c0.clk
		.areset    (),                                                //        areset_conduit.export
		.locked    (),                                                //        locked_conduit.export
		.phasedone ()                                                 //     phasedone_conduit.export
	);

	DECA_QSYS_sw sw (
		.clk        (pll_c1_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_sw_s1_address),     //                  s1.address
		.write_n    (~mm_interconnect_1_sw_s1_write),      //                    .write_n
		.writedata  (mm_interconnect_1_sw_s1_writedata),   //                    .writedata
		.chipselect (mm_interconnect_1_sw_s1_chipselect),  //                    .chipselect
		.readdata   (mm_interconnect_1_sw_s1_readdata),    //                    .readdata
		.in_port    (pio_sw_external_connection_export),   // external_connection.export
		.irq        (irq_synchronizer_001_receiver_irq)    //                 irq.irq
	);

	DECA_QSYS_sysid_qsys sysid_qsys (
		.clock    (pll_c0_clk),                                          //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_qsys_control_slave_address)   //              .address
	);

	DECA_QSYS_timer timer (
		.clk        (pll_c0_clk),                            //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_1_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)               //   irq.irq
	);

	DECA_QSYS_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                        (clk_clk),                                                     //                                      clk_50_clk.clk
		.pll_c0_clk                                            (pll_c0_clk),                                                  //                                          pll_c0.clk
		.jtag_uart_reset_reset_bridge_in_reset_reset           (rst_controller_002_reset_out_reset),                          //           jtag_uart_reset_reset_bridge_in_reset.reset
		.nios2_gen2_reset_reset_bridge_in_reset_reset          (rst_controller_003_reset_out_reset),                          //          nios2_gen2_reset_reset_bridge_in_reset.reset
		.pll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2_gen2_data_master_address                        (nios2_gen2_data_master_address),                              //                          nios2_gen2_data_master.address
		.nios2_gen2_data_master_waitrequest                    (nios2_gen2_data_master_waitrequest),                          //                                                .waitrequest
		.nios2_gen2_data_master_byteenable                     (nios2_gen2_data_master_byteenable),                           //                                                .byteenable
		.nios2_gen2_data_master_read                           (nios2_gen2_data_master_read),                                 //                                                .read
		.nios2_gen2_data_master_readdata                       (nios2_gen2_data_master_readdata),                             //                                                .readdata
		.nios2_gen2_data_master_readdatavalid                  (nios2_gen2_data_master_readdatavalid),                        //                                                .readdatavalid
		.nios2_gen2_data_master_write                          (nios2_gen2_data_master_write),                                //                                                .write
		.nios2_gen2_data_master_writedata                      (nios2_gen2_data_master_writedata),                            //                                                .writedata
		.nios2_gen2_data_master_debugaccess                    (nios2_gen2_data_master_debugaccess),                          //                                                .debugaccess
		.nios2_gen2_instruction_master_address                 (nios2_gen2_instruction_master_address),                       //                   nios2_gen2_instruction_master.address
		.nios2_gen2_instruction_master_waitrequest             (nios2_gen2_instruction_master_waitrequest),                   //                                                .waitrequest
		.nios2_gen2_instruction_master_read                    (nios2_gen2_instruction_master_read),                          //                                                .read
		.nios2_gen2_instruction_master_readdata                (nios2_gen2_instruction_master_readdata),                      //                                                .readdata
		.nios2_gen2_instruction_master_readdatavalid           (nios2_gen2_instruction_master_readdatavalid),                 //                                                .readdatavalid
		.Audio_i2c_avalon_slave_0_address                      (mm_interconnect_0_audio_i2c_avalon_slave_0_address),          //                        Audio_i2c_avalon_slave_0.address
		.Audio_i2c_avalon_slave_0_write                        (mm_interconnect_0_audio_i2c_avalon_slave_0_write),            //                                                .write
		.Audio_i2c_avalon_slave_0_readdata                     (mm_interconnect_0_audio_i2c_avalon_slave_0_readdata),         //                                                .readdata
		.Audio_i2c_avalon_slave_0_writedata                    (mm_interconnect_0_audio_i2c_avalon_slave_0_writedata),        //                                                .writedata
		.Audio_i2c_avalon_slave_0_waitrequest                  (~mm_interconnect_0_audio_i2c_avalon_slave_0_waitrequest),     //                                                .waitrequest
		.Audio_i2c_avalon_slave_0_chipselect                   (mm_interconnect_0_audio_i2c_avalon_slave_0_chipselect),       //                                                .chipselect
		.jtag_uart_avalon_jtag_slave_address                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),       //                     jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),         //                                                .write
		.jtag_uart_avalon_jtag_slave_read                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),          //                                                .read
		.jtag_uart_avalon_jtag_slave_readdata                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),      //                                                .readdata
		.jtag_uart_avalon_jtag_slave_writedata                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),     //                                                .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),   //                                                .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),    //                                                .chipselect
		.mm_clock_crossing_bridge_s0_address                   (mm_interconnect_0_mm_clock_crossing_bridge_s0_address),       //                     mm_clock_crossing_bridge_s0.address
		.mm_clock_crossing_bridge_s0_write                     (mm_interconnect_0_mm_clock_crossing_bridge_s0_write),         //                                                .write
		.mm_clock_crossing_bridge_s0_read                      (mm_interconnect_0_mm_clock_crossing_bridge_s0_read),          //                                                .read
		.mm_clock_crossing_bridge_s0_readdata                  (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata),      //                                                .readdata
		.mm_clock_crossing_bridge_s0_writedata                 (mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata),     //                                                .writedata
		.mm_clock_crossing_bridge_s0_burstcount                (mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount),    //                                                .burstcount
		.mm_clock_crossing_bridge_s0_byteenable                (mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable),    //                                                .byteenable
		.mm_clock_crossing_bridge_s0_readdatavalid             (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid), //                                                .readdatavalid
		.mm_clock_crossing_bridge_s0_waitrequest               (mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest),   //                                                .waitrequest
		.mm_clock_crossing_bridge_s0_debugaccess               (mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess),   //                                                .debugaccess
		.nios2_gen2_debug_mem_slave_address                    (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),        //                      nios2_gen2_debug_mem_slave.address
		.nios2_gen2_debug_mem_slave_write                      (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),          //                                                .write
		.nios2_gen2_debug_mem_slave_read                       (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),           //                                                .read
		.nios2_gen2_debug_mem_slave_readdata                   (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),       //                                                .readdata
		.nios2_gen2_debug_mem_slave_writedata                  (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),      //                                                .writedata
		.nios2_gen2_debug_mem_slave_byteenable                 (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),     //                                                .byteenable
		.nios2_gen2_debug_mem_slave_waitrequest                (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest),    //                                                .waitrequest
		.nios2_gen2_debug_mem_slave_debugaccess                (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess),    //                                                .debugaccess
		.onchip_memory2_s1_address                             (mm_interconnect_0_onchip_memory2_s1_address),                 //                               onchip_memory2_s1.address
		.onchip_memory2_s1_write                               (mm_interconnect_0_onchip_memory2_s1_write),                   //                                                .write
		.onchip_memory2_s1_readdata                            (mm_interconnect_0_onchip_memory2_s1_readdata),                //                                                .readdata
		.onchip_memory2_s1_writedata                           (mm_interconnect_0_onchip_memory2_s1_writedata),               //                                                .writedata
		.onchip_memory2_s1_byteenable                          (mm_interconnect_0_onchip_memory2_s1_byteenable),              //                                                .byteenable
		.onchip_memory2_s1_chipselect                          (mm_interconnect_0_onchip_memory2_s1_chipselect),              //                                                .chipselect
		.onchip_memory2_s1_clken                               (mm_interconnect_0_onchip_memory2_s1_clken),                   //                                                .clken
		.pll_pll_slave_address                                 (mm_interconnect_0_pll_pll_slave_address),                     //                                   pll_pll_slave.address
		.pll_pll_slave_write                                   (mm_interconnect_0_pll_pll_slave_write),                       //                                                .write
		.pll_pll_slave_read                                    (mm_interconnect_0_pll_pll_slave_read),                        //                                                .read
		.pll_pll_slave_readdata                                (mm_interconnect_0_pll_pll_slave_readdata),                    //                                                .readdata
		.pll_pll_slave_writedata                               (mm_interconnect_0_pll_pll_slave_writedata),                   //                                                .writedata
		.pll_audio_pll_slave_address                           (mm_interconnect_0_pll_audio_pll_slave_address),               //                             pll_audio_pll_slave.address
		.pll_audio_pll_slave_write                             (mm_interconnect_0_pll_audio_pll_slave_write),                 //                                                .write
		.pll_audio_pll_slave_read                              (mm_interconnect_0_pll_audio_pll_slave_read),                  //                                                .read
		.pll_audio_pll_slave_readdata                          (mm_interconnect_0_pll_audio_pll_slave_readdata),              //                                                .readdata
		.pll_audio_pll_slave_writedata                         (mm_interconnect_0_pll_audio_pll_slave_writedata)              //                                                .writedata
	);

	DECA_QSYS_mm_interconnect_1 mm_interconnect_1 (
		.pll_c0_clk                                                    (pll_c0_clk),                                          //                                                  pll_c0.clk
		.pll_c1_clk                                                    (pll_c1_clk),                                          //                                                  pll_c1.clk
		.mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                  // mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset.reset
		.sysid_qsys_reset_reset_bridge_in_reset_reset                  (rst_controller_002_reset_out_reset),                  //                  sysid_qsys_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_m0_address                           (mm_clock_crossing_bridge_m0_address),                 //                             mm_clock_crossing_bridge_m0.address
		.mm_clock_crossing_bridge_m0_waitrequest                       (mm_clock_crossing_bridge_m0_waitrequest),             //                                                        .waitrequest
		.mm_clock_crossing_bridge_m0_burstcount                        (mm_clock_crossing_bridge_m0_burstcount),              //                                                        .burstcount
		.mm_clock_crossing_bridge_m0_byteenable                        (mm_clock_crossing_bridge_m0_byteenable),              //                                                        .byteenable
		.mm_clock_crossing_bridge_m0_read                              (mm_clock_crossing_bridge_m0_read),                    //                                                        .read
		.mm_clock_crossing_bridge_m0_readdata                          (mm_clock_crossing_bridge_m0_readdata),                //                                                        .readdata
		.mm_clock_crossing_bridge_m0_readdatavalid                     (mm_clock_crossing_bridge_m0_readdatavalid),           //                                                        .readdatavalid
		.mm_clock_crossing_bridge_m0_write                             (mm_clock_crossing_bridge_m0_write),                   //                                                        .write
		.mm_clock_crossing_bridge_m0_writedata                         (mm_clock_crossing_bridge_m0_writedata),               //                                                        .writedata
		.mm_clock_crossing_bridge_m0_debugaccess                       (mm_clock_crossing_bridge_m0_debugaccess),             //                                                        .debugaccess
		.audio_reset_n_s1_address                                      (mm_interconnect_1_audio_reset_n_s1_address),          //                                        audio_reset_n_s1.address
		.audio_reset_n_s1_write                                        (mm_interconnect_1_audio_reset_n_s1_write),            //                                                        .write
		.audio_reset_n_s1_readdata                                     (mm_interconnect_1_audio_reset_n_s1_readdata),         //                                                        .readdata
		.audio_reset_n_s1_writedata                                    (mm_interconnect_1_audio_reset_n_s1_writedata),        //                                                        .writedata
		.audio_reset_n_s1_chipselect                                   (mm_interconnect_1_audio_reset_n_s1_chipselect),       //                                                        .chipselect
		.key_s1_address                                                (mm_interconnect_1_key_s1_address),                    //                                                  key_s1.address
		.key_s1_write                                                  (mm_interconnect_1_key_s1_write),                      //                                                        .write
		.key_s1_readdata                                               (mm_interconnect_1_key_s1_readdata),                   //                                                        .readdata
		.key_s1_writedata                                              (mm_interconnect_1_key_s1_writedata),                  //                                                        .writedata
		.key_s1_chipselect                                             (mm_interconnect_1_key_s1_chipselect),                 //                                                        .chipselect
		.led_s1_address                                                (mm_interconnect_1_led_s1_address),                    //                                                  led_s1.address
		.led_s1_write                                                  (mm_interconnect_1_led_s1_write),                      //                                                        .write
		.led_s1_readdata                                               (mm_interconnect_1_led_s1_readdata),                   //                                                        .readdata
		.led_s1_writedata                                              (mm_interconnect_1_led_s1_writedata),                  //                                                        .writedata
		.led_s1_chipselect                                             (mm_interconnect_1_led_s1_chipselect),                 //                                                        .chipselect
		.sw_s1_address                                                 (mm_interconnect_1_sw_s1_address),                     //                                                   sw_s1.address
		.sw_s1_write                                                   (mm_interconnect_1_sw_s1_write),                       //                                                        .write
		.sw_s1_readdata                                                (mm_interconnect_1_sw_s1_readdata),                    //                                                        .readdata
		.sw_s1_writedata                                               (mm_interconnect_1_sw_s1_writedata),                   //                                                        .writedata
		.sw_s1_chipselect                                              (mm_interconnect_1_sw_s1_chipselect),                  //                                                        .chipselect
		.sysid_qsys_control_slave_address                              (mm_interconnect_1_sysid_qsys_control_slave_address),  //                                sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                             (mm_interconnect_1_sysid_qsys_control_slave_readdata), //                                                        .readdata
		.timer_s1_address                                              (mm_interconnect_1_timer_s1_address),                  //                                                timer_s1.address
		.timer_s1_write                                                (mm_interconnect_1_timer_s1_write),                    //                                                        .write
		.timer_s1_readdata                                             (mm_interconnect_1_timer_s1_readdata),                 //                                                        .readdata
		.timer_s1_writedata                                            (mm_interconnect_1_timer_s1_writedata),                //                                                        .writedata
		.timer_s1_chipselect                                           (mm_interconnect_1_timer_s1_chipselect)                //                                                        .chipselect
	);

	DECA_QSYS_irq_mapper irq_mapper (
		.clk           (pll_c0_clk),                         //       clk.clk
		.reset         (rst_controller_003_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (nios2_gen2_irq_irq)                  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (pll_c0_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_003_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (pll_c1_clk),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_003_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (pll_c1_clk),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_003_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_c1_clk),                         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (pll_c0_clk),                             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset),   // reset_in1.reset
		.clk            (pll_c0_clk),                             //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_003_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
