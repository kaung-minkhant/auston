// deca_qsys.v

// Generated using ACDS version 15.0 143

`timescale 1 ps / 1 ps
module deca_qsys (
		input  wire        clk_clk,                                       //                             clk.clk
		input  wire [3:0]  ddr3_status_external_connection_export,        // ddr3_status_external_connection.export
		input  wire [1:0]  key_external_connection_export,                //         key_external_connection.export
		input  wire        mem_if_ddr3_emif_pll_ref_clk_clk,              //    mem_if_ddr3_emif_pll_ref_clk.clk
		output wire        mem_if_ddr3_emif_pll_sharing_pll_mem_clk,      //    mem_if_ddr3_emif_pll_sharing.pll_mem_clk
		output wire        mem_if_ddr3_emif_pll_sharing_pll_write_clk,    //                                .pll_write_clk
		output wire        mem_if_ddr3_emif_pll_sharing_pll_locked,       //                                .pll_locked
		output wire        mem_if_ddr3_emif_pll_sharing_pll_capture0_clk, //                                .pll_capture0_clk
		output wire        mem_if_ddr3_emif_pll_sharing_pll_capture1_clk, //                                .pll_capture1_clk
		output wire        mem_if_ddr3_emif_status_local_init_done,       //         mem_if_ddr3_emif_status.local_init_done
		output wire        mem_if_ddr3_emif_status_local_cal_success,     //                                .local_cal_success
		output wire        mem_if_ddr3_emif_status_local_cal_fail,        //                                .local_cal_fail
		output wire [14:0] memory_mem_a,                                  //                          memory.mem_a
		output wire [2:0]  memory_mem_ba,                                 //                                .mem_ba
		inout  wire [0:0]  memory_mem_ck,                                 //                                .mem_ck
		inout  wire [0:0]  memory_mem_ck_n,                               //                                .mem_ck_n
		output wire [0:0]  memory_mem_cke,                                //                                .mem_cke
		output wire [0:0]  memory_mem_cs_n,                               //                                .mem_cs_n
		output wire [1:0]  memory_mem_dm,                                 //                                .mem_dm
		output wire [0:0]  memory_mem_ras_n,                              //                                .mem_ras_n
		output wire [0:0]  memory_mem_cas_n,                              //                                .mem_cas_n
		output wire [0:0]  memory_mem_we_n,                               //                                .mem_we_n
		output wire        memory_mem_reset_n,                            //                                .mem_reset_n
		inout  wire [15:0] memory_mem_dq,                                 //                                .mem_dq
		inout  wire [1:0]  memory_mem_dqs,                                //                                .mem_dqs
		inout  wire [1:0]  memory_mem_dqs_n,                              //                                .mem_dqs_n
		output wire [0:0]  memory_mem_odt,                                //                                .mem_odt
		input  wire        reset_reset_n                                  //                           reset.reset_n
	);

	wire         mem_if_ddr3_emif_afi_half_clk_clk;                                // mem_if_ddr3_emif:afi_half_clk -> [mm_clock_crossing_bridge_ddr3:m0_clk, rst_controller_002:clk]
	wire         altpll_sys_c0_clk;                                                // altpll_sys:c0 -> [irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, mm_clock_crossing_bridge_ddr3:s0_clk, mm_clock_crossing_bridge_io:s0_clk, mm_interconnect_0:altpll_sys_c0_clk, nios2_gen2:clk, onchip_memory2:clk, rst_controller_003:clk, rst_controller_004:clk]
	wire         altpll_sys_c1_clk;                                                // altpll_sys:c1 -> [ddr3_status:clk, irq_synchronizer_001:receiver_clk, jtag_uart:clk, key:clk, mm_clock_crossing_bridge_io:m0_clk, mm_interconnect_1:altpll_sys_c1_clk, rst_controller_001:clk, sysid_qsys:clock]
	wire  [31:0] nios2_gen2_data_master_readdata;                                  // mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	wire         nios2_gen2_data_master_waitrequest;                               // mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	wire         nios2_gen2_data_master_debugaccess;                               // nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
	wire  [29:0] nios2_gen2_data_master_address;                                   // nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
	wire   [3:0] nios2_gen2_data_master_byteenable;                                // nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
	wire         nios2_gen2_data_master_read;                                      // nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
	wire         nios2_gen2_data_master_readdatavalid;                             // mm_interconnect_0:nios2_gen2_data_master_readdatavalid -> nios2_gen2:d_readdatavalid
	wire         nios2_gen2_data_master_write;                                     // nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
	wire  [31:0] nios2_gen2_data_master_writedata;                                 // nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
	wire  [31:0] nios2_gen2_instruction_master_readdata;                           // mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	wire         nios2_gen2_instruction_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	wire  [29:0] nios2_gen2_instruction_master_address;                            // nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
	wire         nios2_gen2_instruction_master_read;                               // nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
	wire         nios2_gen2_instruction_master_readdatavalid;                      // mm_interconnect_0:nios2_gen2_instruction_master_readdatavalid -> nios2_gen2:i_readdatavalid
	wire         mm_interconnect_0_mem_if_ddr3_emif_avl_beginbursttransfer;        // mm_interconnect_0:mem_if_ddr3_emif_avl_beginbursttransfer -> mem_if_ddr3_emif:avl_burstbegin
	wire  [63:0] mm_interconnect_0_mem_if_ddr3_emif_avl_readdata;                  // mem_if_ddr3_emif:avl_rdata -> mm_interconnect_0:mem_if_ddr3_emif_avl_readdata
	wire         mm_interconnect_0_mem_if_ddr3_emif_avl_waitrequest;               // mem_if_ddr3_emif:avl_ready -> mm_interconnect_0:mem_if_ddr3_emif_avl_waitrequest
	wire  [25:0] mm_interconnect_0_mem_if_ddr3_emif_avl_address;                   // mm_interconnect_0:mem_if_ddr3_emif_avl_address -> mem_if_ddr3_emif:avl_addr
	wire         mm_interconnect_0_mem_if_ddr3_emif_avl_read;                      // mm_interconnect_0:mem_if_ddr3_emif_avl_read -> mem_if_ddr3_emif:avl_read_req
	wire   [7:0] mm_interconnect_0_mem_if_ddr3_emif_avl_byteenable;                // mm_interconnect_0:mem_if_ddr3_emif_avl_byteenable -> mem_if_ddr3_emif:avl_be
	wire         mm_interconnect_0_mem_if_ddr3_emif_avl_readdatavalid;             // mem_if_ddr3_emif:avl_rdata_valid -> mm_interconnect_0:mem_if_ddr3_emif_avl_readdatavalid
	wire         mm_interconnect_0_mem_if_ddr3_emif_avl_write;                     // mm_interconnect_0:mem_if_ddr3_emif_avl_write -> mem_if_ddr3_emif:avl_write_req
	wire  [63:0] mm_interconnect_0_mem_if_ddr3_emif_avl_writedata;                 // mm_interconnect_0:mem_if_ddr3_emif_avl_writedata -> mem_if_ddr3_emif:avl_wdata
	wire   [2:0] mm_interconnect_0_mem_if_ddr3_emif_avl_burstcount;                // mm_interconnect_0:mem_if_ddr3_emif_avl_burstcount -> mem_if_ddr3_emif:avl_size
	wire         mem_if_ddr3_emif_afi_clk_clk;                                     // mem_if_ddr3_emif:afi_clk -> [mm_interconnect_0:mem_if_ddr3_emif_afi_clk_clk, rst_controller_005:clk]
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata;            // nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest;         // nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess;         // mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_address;             // mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_read;                // mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable;          // mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_write;               // mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata;           // mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_sys_pll_slave_readdata;                  // altpll_sys:readdata -> mm_interconnect_0:altpll_sys_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_sys_pll_slave_address;                   // mm_interconnect_0:altpll_sys_pll_slave_address -> altpll_sys:address
	wire         mm_interconnect_0_altpll_sys_pll_slave_read;                      // mm_interconnect_0:altpll_sys_pll_slave_read -> altpll_sys:read
	wire         mm_interconnect_0_altpll_sys_pll_slave_write;                     // mm_interconnect_0:altpll_sys_pll_slave_write -> altpll_sys:write
	wire  [31:0] mm_interconnect_0_altpll_sys_pll_slave_writedata;                 // mm_interconnect_0:altpll_sys_pll_slave_writedata -> altpll_sys:writedata
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_readdata;      // mm_clock_crossing_bridge_ddr3:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_ddr3_s0_readdata
	wire         mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_waitrequest;   // mm_clock_crossing_bridge_ddr3:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_ddr3_s0_waitrequest
	wire         mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_debugaccess;   // mm_interconnect_0:mm_clock_crossing_bridge_ddr3_s0_debugaccess -> mm_clock_crossing_bridge_ddr3:s0_debugaccess
	wire   [9:0] mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_address;       // mm_interconnect_0:mm_clock_crossing_bridge_ddr3_s0_address -> mm_clock_crossing_bridge_ddr3:s0_address
	wire         mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_read;          // mm_interconnect_0:mm_clock_crossing_bridge_ddr3_s0_read -> mm_clock_crossing_bridge_ddr3:s0_read
	wire   [3:0] mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_byteenable;    // mm_interconnect_0:mm_clock_crossing_bridge_ddr3_s0_byteenable -> mm_clock_crossing_bridge_ddr3:s0_byteenable
	wire         mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_readdatavalid; // mm_clock_crossing_bridge_ddr3:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_ddr3_s0_readdatavalid
	wire         mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_write;         // mm_interconnect_0:mm_clock_crossing_bridge_ddr3_s0_write -> mm_clock_crossing_bridge_ddr3:s0_write
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_writedata;     // mm_interconnect_0:mm_clock_crossing_bridge_ddr3_s0_writedata -> mm_clock_crossing_bridge_ddr3:s0_writedata
	wire   [0:0] mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_burstcount;    // mm_interconnect_0:mm_clock_crossing_bridge_ddr3_s0_burstcount -> mm_clock_crossing_bridge_ddr3:s0_burstcount
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_io_s0_readdata;        // mm_clock_crossing_bridge_io:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_io_s0_readdata
	wire         mm_interconnect_0_mm_clock_crossing_bridge_io_s0_waitrequest;     // mm_clock_crossing_bridge_io:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_io_s0_waitrequest
	wire         mm_interconnect_0_mm_clock_crossing_bridge_io_s0_debugaccess;     // mm_interconnect_0:mm_clock_crossing_bridge_io_s0_debugaccess -> mm_clock_crossing_bridge_io:s0_debugaccess
	wire   [9:0] mm_interconnect_0_mm_clock_crossing_bridge_io_s0_address;         // mm_interconnect_0:mm_clock_crossing_bridge_io_s0_address -> mm_clock_crossing_bridge_io:s0_address
	wire         mm_interconnect_0_mm_clock_crossing_bridge_io_s0_read;            // mm_interconnect_0:mm_clock_crossing_bridge_io_s0_read -> mm_clock_crossing_bridge_io:s0_read
	wire   [3:0] mm_interconnect_0_mm_clock_crossing_bridge_io_s0_byteenable;      // mm_interconnect_0:mm_clock_crossing_bridge_io_s0_byteenable -> mm_clock_crossing_bridge_io:s0_byteenable
	wire         mm_interconnect_0_mm_clock_crossing_bridge_io_s0_readdatavalid;   // mm_clock_crossing_bridge_io:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_io_s0_readdatavalid
	wire         mm_interconnect_0_mm_clock_crossing_bridge_io_s0_write;           // mm_interconnect_0:mm_clock_crossing_bridge_io_s0_write -> mm_clock_crossing_bridge_io:s0_write
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_io_s0_writedata;       // mm_interconnect_0:mm_clock_crossing_bridge_io_s0_writedata -> mm_clock_crossing_bridge_io:s0_writedata
	wire   [0:0] mm_interconnect_0_mm_clock_crossing_bridge_io_s0_burstcount;      // mm_interconnect_0:mm_clock_crossing_bridge_io_s0_burstcount -> mm_clock_crossing_bridge_io:s0_burstcount
	wire         mm_interconnect_0_onchip_memory2_s1_chipselect;                   // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;                     // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire  [14:0] mm_interconnect_0_onchip_memory2_s1_address;                      // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;                   // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire         mm_interconnect_0_onchip_memory2_s1_write;                        // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;                    // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire         mm_interconnect_0_onchip_memory2_s1_clken;                        // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire         mm_clock_crossing_bridge_io_m0_waitrequest;                       // mm_interconnect_1:mm_clock_crossing_bridge_io_m0_waitrequest -> mm_clock_crossing_bridge_io:m0_waitrequest
	wire  [31:0] mm_clock_crossing_bridge_io_m0_readdata;                          // mm_interconnect_1:mm_clock_crossing_bridge_io_m0_readdata -> mm_clock_crossing_bridge_io:m0_readdata
	wire         mm_clock_crossing_bridge_io_m0_debugaccess;                       // mm_clock_crossing_bridge_io:m0_debugaccess -> mm_interconnect_1:mm_clock_crossing_bridge_io_m0_debugaccess
	wire   [9:0] mm_clock_crossing_bridge_io_m0_address;                           // mm_clock_crossing_bridge_io:m0_address -> mm_interconnect_1:mm_clock_crossing_bridge_io_m0_address
	wire         mm_clock_crossing_bridge_io_m0_read;                              // mm_clock_crossing_bridge_io:m0_read -> mm_interconnect_1:mm_clock_crossing_bridge_io_m0_read
	wire   [3:0] mm_clock_crossing_bridge_io_m0_byteenable;                        // mm_clock_crossing_bridge_io:m0_byteenable -> mm_interconnect_1:mm_clock_crossing_bridge_io_m0_byteenable
	wire         mm_clock_crossing_bridge_io_m0_readdatavalid;                     // mm_interconnect_1:mm_clock_crossing_bridge_io_m0_readdatavalid -> mm_clock_crossing_bridge_io:m0_readdatavalid
	wire  [31:0] mm_clock_crossing_bridge_io_m0_writedata;                         // mm_clock_crossing_bridge_io:m0_writedata -> mm_interconnect_1:mm_clock_crossing_bridge_io_m0_writedata
	wire         mm_clock_crossing_bridge_io_m0_write;                             // mm_clock_crossing_bridge_io:m0_write -> mm_interconnect_1:mm_clock_crossing_bridge_io_m0_write
	wire   [0:0] mm_clock_crossing_bridge_io_m0_burstcount;                        // mm_clock_crossing_bridge_io:m0_burstcount -> mm_interconnect_1:mm_clock_crossing_bridge_io_m0_burstcount
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;         // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;           // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest;        // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;            // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;               // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;              // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;          // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_1_sysid_qsys_control_slave_readdata;              // sysid_qsys:readdata -> mm_interconnect_1:sysid_qsys_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_qsys_control_slave_address;               // mm_interconnect_1:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire         mm_interconnect_1_timer_s1_chipselect;                            // mm_interconnect_1:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_1_timer_s1_readdata;                              // timer:readdata -> mm_interconnect_1:timer_s1_readdata
	wire   [2:0] mm_interconnect_1_timer_s1_address;                               // mm_interconnect_1:timer_s1_address -> timer:address
	wire         mm_interconnect_1_timer_s1_write;                                 // mm_interconnect_1:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_1_timer_s1_writedata;                             // mm_interconnect_1:timer_s1_writedata -> timer:writedata
	wire  [31:0] mm_interconnect_1_key_s1_readdata;                                // key:readdata -> mm_interconnect_1:key_s1_readdata
	wire   [1:0] mm_interconnect_1_key_s1_address;                                 // mm_interconnect_1:key_s1_address -> key:address
	wire  [31:0] mm_interconnect_1_ddr3_status_s1_readdata;                        // ddr3_status:readdata -> mm_interconnect_1:ddr3_status_s1_readdata
	wire   [1:0] mm_interconnect_1_ddr3_status_s1_address;                         // mm_interconnect_1:ddr3_status_s1_address -> ddr3_status:address
	wire  [31:0] nios2_gen2_irq_irq;                                               // irq_mapper:sender_irq -> nios2_gen2:irq
	wire         irq_mapper_receiver0_irq;                                         // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                    // timer:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver1_irq;                                         // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                // jtag_uart:av_irq -> irq_synchronizer_001:receiver_irq
	wire         rst_controller_reset_out_reset;                                   // rst_controller:reset_out -> [altpll_sys:reset, irq_synchronizer:receiver_reset, mm_interconnect_0:altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset, mm_interconnect_1:timer_reset_reset_bridge_in_reset_reset, timer:reset_n]
	wire         rst_controller_001_reset_out_reset;                               // rst_controller_001:reset_out -> [ddr3_status:reset_n, irq_synchronizer_001:receiver_reset, jtag_uart:rst_n, key:reset_n, mm_clock_crossing_bridge_io:m0_reset, mm_interconnect_1:mm_clock_crossing_bridge_io_m0_reset_reset_bridge_in_reset_reset, sysid_qsys:reset_n]
	wire         rst_controller_002_reset_out_reset;                               // rst_controller_002:reset_out -> mm_clock_crossing_bridge_ddr3:m0_reset
	wire         rst_controller_003_reset_out_reset;                               // rst_controller_003:reset_out -> [mm_clock_crossing_bridge_ddr3:s0_reset, mm_clock_crossing_bridge_io:s0_reset, mm_interconnect_0:mm_clock_crossing_bridge_ddr3_s0_reset_reset_bridge_in_reset_reset, onchip_memory2:reset, rst_translator:in_reset]
	wire         rst_controller_003_reset_out_reset_req;                           // rst_controller_003:reset_req -> [onchip_memory2:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_004_reset_out_reset;                               // rst_controller_004:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_interconnect_0:nios2_gen2_reset_reset_bridge_in_reset_reset, nios2_gen2:reset_n, rst_translator_001:in_reset]
	wire         rst_controller_004_reset_out_reset_req;                           // rst_controller_004:reset_req -> [nios2_gen2:reset_req, rst_translator_001:reset_req_in]
	wire         nios2_gen2_debug_reset_request_reset;                             // nios2_gen2:debug_reset_request -> rst_controller_004:reset_in1
	wire         rst_controller_005_reset_out_reset;                               // rst_controller_005:reset_out -> [mm_interconnect_0:mem_if_ddr3_emif_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mem_if_ddr3_emif_soft_reset_reset_bridge_in_reset_reset]

	deca_qsys_altpll_sys altpll_sys (
		.clk       (clk_clk),                                          //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),                   // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_sys_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_sys_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_sys_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_sys_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_sys_pll_slave_writedata), //                      .writedata
		.c0        (altpll_sys_c0_clk),                                //                    c0.clk
		.c1        (altpll_sys_c1_clk),                                //                    c1.clk
		.areset    (),                                                 //        areset_conduit.export
		.locked    (),                                                 //        locked_conduit.export
		.phasedone ()                                                  //     phasedone_conduit.export
	);

	deca_qsys_ddr3_status ddr3_status (
		.clk      (altpll_sys_c1_clk),                         //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_1_ddr3_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_ddr3_status_s1_readdata), //                    .readdata
		.in_port  (ddr3_status_external_connection_export)     // external_connection.export
	);

	deca_qsys_jtag_uart jtag_uart (
		.clk            (altpll_sys_c1_clk),                                         //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_001_receiver_irq)                          //               irq.irq
	);

	deca_qsys_key key (
		.clk      (altpll_sys_c1_clk),                   //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_1_key_s1_address),    //                  s1.address
		.readdata (mm_interconnect_1_key_s1_readdata),   //                    .readdata
		.in_port  (key_external_connection_export)       // external_connection.export
	);

	deca_qsys_mem_if_ddr3_emif mem_if_ddr3_emif (
		.pll_ref_clk        (mem_if_ddr3_emif_pll_ref_clk_clk),                          //      pll_ref_clk.clk
		.global_reset_n     (reset_reset_n),                                             //     global_reset.reset_n
		.soft_reset_n       (reset_reset_n),                                             //       soft_reset.reset_n
		.afi_clk            (mem_if_ddr3_emif_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk       (mem_if_ddr3_emif_afi_half_clk_clk),                         //     afi_half_clk.clk
		.afi_reset_n        (),                                                          //        afi_reset.reset_n
		.afi_reset_export_n (),                                                          // afi_reset_export.reset_n
		.mem_a              (memory_mem_a),                                              //           memory.mem_a
		.mem_ba             (memory_mem_ba),                                             //                 .mem_ba
		.mem_ck             (memory_mem_ck),                                             //                 .mem_ck
		.mem_ck_n           (memory_mem_ck_n),                                           //                 .mem_ck_n
		.mem_cke            (memory_mem_cke),                                            //                 .mem_cke
		.mem_cs_n           (memory_mem_cs_n),                                           //                 .mem_cs_n
		.mem_dm             (memory_mem_dm),                                             //                 .mem_dm
		.mem_ras_n          (memory_mem_ras_n),                                          //                 .mem_ras_n
		.mem_cas_n          (memory_mem_cas_n),                                          //                 .mem_cas_n
		.mem_we_n           (memory_mem_we_n),                                           //                 .mem_we_n
		.mem_reset_n        (memory_mem_reset_n),                                        //                 .mem_reset_n
		.mem_dq             (memory_mem_dq),                                             //                 .mem_dq
		.mem_dqs            (memory_mem_dqs),                                            //                 .mem_dqs
		.mem_dqs_n          (memory_mem_dqs_n),                                          //                 .mem_dqs_n
		.mem_odt            (memory_mem_odt),                                            //                 .mem_odt
		.avl_ready          (mm_interconnect_0_mem_if_ddr3_emif_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin     (mm_interconnect_0_mem_if_ddr3_emif_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr           (mm_interconnect_0_mem_if_ddr3_emif_avl_address),            //                 .address
		.avl_rdata_valid    (mm_interconnect_0_mem_if_ddr3_emif_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata          (mm_interconnect_0_mem_if_ddr3_emif_avl_readdata),           //                 .readdata
		.avl_wdata          (mm_interconnect_0_mem_if_ddr3_emif_avl_writedata),          //                 .writedata
		.avl_be             (mm_interconnect_0_mem_if_ddr3_emif_avl_byteenable),         //                 .byteenable
		.avl_read_req       (mm_interconnect_0_mem_if_ddr3_emif_avl_read),               //                 .read
		.avl_write_req      (mm_interconnect_0_mem_if_ddr3_emif_avl_write),              //                 .write
		.avl_size           (mm_interconnect_0_mem_if_ddr3_emif_avl_burstcount),         //                 .burstcount
		.local_init_done    (mem_if_ddr3_emif_status_local_init_done),                   //           status.local_init_done
		.local_cal_success  (mem_if_ddr3_emif_status_local_cal_success),                 //                 .local_cal_success
		.local_cal_fail     (mem_if_ddr3_emif_status_local_cal_fail),                    //                 .local_cal_fail
		.pll_mem_clk        (mem_if_ddr3_emif_pll_sharing_pll_mem_clk),                  //      pll_sharing.pll_mem_clk
		.pll_write_clk      (mem_if_ddr3_emif_pll_sharing_pll_write_clk),                //                 .pll_write_clk
		.pll_locked         (mem_if_ddr3_emif_pll_sharing_pll_locked),                   //                 .pll_locked
		.pll_capture0_clk   (mem_if_ddr3_emif_pll_sharing_pll_capture0_clk),             //                 .pll_capture0_clk
		.pll_capture1_clk   (mem_if_ddr3_emif_pll_sharing_pll_capture1_clk)              //                 .pll_capture1_clk
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge_ddr3 (
		.m0_clk           (mem_if_ddr3_emif_afi_half_clk_clk),                                //   m0_clk.clk
		.m0_reset         (rst_controller_002_reset_out_reset),                               // m0_reset.reset
		.s0_clk           (altpll_sys_c0_clk),                                                //   s0_clk.clk
		.s0_reset         (rst_controller_003_reset_out_reset),                               // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (),                                                                 //       m0.waitrequest
		.m0_readdata      (),                                                                 //         .readdata
		.m0_readdatavalid (),                                                                 //         .readdatavalid
		.m0_burstcount    (),                                                                 //         .burstcount
		.m0_writedata     (),                                                                 //         .writedata
		.m0_address       (),                                                                 //         .address
		.m0_write         (),                                                                 //         .write
		.m0_read          (),                                                                 //         .read
		.m0_byteenable    (),                                                                 //         .byteenable
		.m0_debugaccess   ()                                                                  //         .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge_io (
		.m0_clk           (altpll_sys_c1_clk),                                              //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                             // m0_reset.reset
		.s0_clk           (altpll_sys_c0_clk),                                              //   s0_clk.clk
		.s0_reset         (rst_controller_003_reset_out_reset),                             // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_io_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_io_m0_readdata),                        //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_io_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_io_m0_burstcount),                      //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_io_m0_writedata),                       //         .writedata
		.m0_address       (mm_clock_crossing_bridge_io_m0_address),                         //         .address
		.m0_write         (mm_clock_crossing_bridge_io_m0_write),                           //         .write
		.m0_read          (mm_clock_crossing_bridge_io_m0_read),                            //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_io_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_io_m0_debugaccess)                      //         .debugaccess
	);

	deca_qsys_nios2_gen2 nios2_gen2 (
		.clk                                 (altpll_sys_c0_clk),                                        //                       clk.clk
		.reset_n                             (~rst_controller_004_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_004_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_gen2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	deca_qsys_onchip_memory2 onchip_memory2 (
		.clk        (altpll_sys_c0_clk),                              //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_003_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_003_reset_out_reset_req)          //       .reset_req
	);

	deca_qsys_sysid_qsys sysid_qsys (
		.clock    (altpll_sys_c1_clk),                                   //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_qsys_control_slave_address)   //              .address
	);

	deca_qsys_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_1_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)          //   irq.irq
	);

	deca_qsys_mm_interconnect_0 mm_interconnect_0 (
		.altpll_sys_c0_clk                                                  (altpll_sys_c0_clk),                                                //                                                altpll_sys_c0.clk
		.clk_50_clk_clk                                                     (clk_clk),                                                          //                                                   clk_50_clk.clk
		.mem_if_ddr3_emif_afi_clk_clk                                       (mem_if_ddr3_emif_afi_clk_clk),                                     //                                     mem_if_ddr3_emif_afi_clk.clk
		.altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                                   //       altpll_sys_inclk_interface_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_avl_translator_reset_reset_bridge_in_reset_reset  (rst_controller_005_reset_out_reset),                               //  mem_if_ddr3_emif_avl_translator_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_soft_reset_reset_bridge_in_reset_reset            (rst_controller_005_reset_out_reset),                               //            mem_if_ddr3_emif_soft_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_ddr3_s0_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),                               // mm_clock_crossing_bridge_ddr3_s0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_reset_reset_bridge_in_reset_reset                       (rst_controller_004_reset_out_reset),                               //                       nios2_gen2_reset_reset_bridge_in_reset.reset
		.nios2_gen2_data_master_address                                     (nios2_gen2_data_master_address),                                   //                                       nios2_gen2_data_master.address
		.nios2_gen2_data_master_waitrequest                                 (nios2_gen2_data_master_waitrequest),                               //                                                             .waitrequest
		.nios2_gen2_data_master_byteenable                                  (nios2_gen2_data_master_byteenable),                                //                                                             .byteenable
		.nios2_gen2_data_master_read                                        (nios2_gen2_data_master_read),                                      //                                                             .read
		.nios2_gen2_data_master_readdata                                    (nios2_gen2_data_master_readdata),                                  //                                                             .readdata
		.nios2_gen2_data_master_readdatavalid                               (nios2_gen2_data_master_readdatavalid),                             //                                                             .readdatavalid
		.nios2_gen2_data_master_write                                       (nios2_gen2_data_master_write),                                     //                                                             .write
		.nios2_gen2_data_master_writedata                                   (nios2_gen2_data_master_writedata),                                 //                                                             .writedata
		.nios2_gen2_data_master_debugaccess                                 (nios2_gen2_data_master_debugaccess),                               //                                                             .debugaccess
		.nios2_gen2_instruction_master_address                              (nios2_gen2_instruction_master_address),                            //                                nios2_gen2_instruction_master.address
		.nios2_gen2_instruction_master_waitrequest                          (nios2_gen2_instruction_master_waitrequest),                        //                                                             .waitrequest
		.nios2_gen2_instruction_master_read                                 (nios2_gen2_instruction_master_read),                               //                                                             .read
		.nios2_gen2_instruction_master_readdata                             (nios2_gen2_instruction_master_readdata),                           //                                                             .readdata
		.nios2_gen2_instruction_master_readdatavalid                        (nios2_gen2_instruction_master_readdatavalid),                      //                                                             .readdatavalid
		.altpll_sys_pll_slave_address                                       (mm_interconnect_0_altpll_sys_pll_slave_address),                   //                                         altpll_sys_pll_slave.address
		.altpll_sys_pll_slave_write                                         (mm_interconnect_0_altpll_sys_pll_slave_write),                     //                                                             .write
		.altpll_sys_pll_slave_read                                          (mm_interconnect_0_altpll_sys_pll_slave_read),                      //                                                             .read
		.altpll_sys_pll_slave_readdata                                      (mm_interconnect_0_altpll_sys_pll_slave_readdata),                  //                                                             .readdata
		.altpll_sys_pll_slave_writedata                                     (mm_interconnect_0_altpll_sys_pll_slave_writedata),                 //                                                             .writedata
		.mem_if_ddr3_emif_avl_address                                       (mm_interconnect_0_mem_if_ddr3_emif_avl_address),                   //                                         mem_if_ddr3_emif_avl.address
		.mem_if_ddr3_emif_avl_write                                         (mm_interconnect_0_mem_if_ddr3_emif_avl_write),                     //                                                             .write
		.mem_if_ddr3_emif_avl_read                                          (mm_interconnect_0_mem_if_ddr3_emif_avl_read),                      //                                                             .read
		.mem_if_ddr3_emif_avl_readdata                                      (mm_interconnect_0_mem_if_ddr3_emif_avl_readdata),                  //                                                             .readdata
		.mem_if_ddr3_emif_avl_writedata                                     (mm_interconnect_0_mem_if_ddr3_emif_avl_writedata),                 //                                                             .writedata
		.mem_if_ddr3_emif_avl_beginbursttransfer                            (mm_interconnect_0_mem_if_ddr3_emif_avl_beginbursttransfer),        //                                                             .beginbursttransfer
		.mem_if_ddr3_emif_avl_burstcount                                    (mm_interconnect_0_mem_if_ddr3_emif_avl_burstcount),                //                                                             .burstcount
		.mem_if_ddr3_emif_avl_byteenable                                    (mm_interconnect_0_mem_if_ddr3_emif_avl_byteenable),                //                                                             .byteenable
		.mem_if_ddr3_emif_avl_readdatavalid                                 (mm_interconnect_0_mem_if_ddr3_emif_avl_readdatavalid),             //                                                             .readdatavalid
		.mem_if_ddr3_emif_avl_waitrequest                                   (~mm_interconnect_0_mem_if_ddr3_emif_avl_waitrequest),              //                                                             .waitrequest
		.mm_clock_crossing_bridge_ddr3_s0_address                           (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_address),       //                             mm_clock_crossing_bridge_ddr3_s0.address
		.mm_clock_crossing_bridge_ddr3_s0_write                             (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_write),         //                                                             .write
		.mm_clock_crossing_bridge_ddr3_s0_read                              (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_read),          //                                                             .read
		.mm_clock_crossing_bridge_ddr3_s0_readdata                          (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_readdata),      //                                                             .readdata
		.mm_clock_crossing_bridge_ddr3_s0_writedata                         (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_writedata),     //                                                             .writedata
		.mm_clock_crossing_bridge_ddr3_s0_burstcount                        (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_burstcount),    //                                                             .burstcount
		.mm_clock_crossing_bridge_ddr3_s0_byteenable                        (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_byteenable),    //                                                             .byteenable
		.mm_clock_crossing_bridge_ddr3_s0_readdatavalid                     (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_readdatavalid), //                                                             .readdatavalid
		.mm_clock_crossing_bridge_ddr3_s0_waitrequest                       (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_waitrequest),   //                                                             .waitrequest
		.mm_clock_crossing_bridge_ddr3_s0_debugaccess                       (mm_interconnect_0_mm_clock_crossing_bridge_ddr3_s0_debugaccess),   //                                                             .debugaccess
		.mm_clock_crossing_bridge_io_s0_address                             (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_address),         //                               mm_clock_crossing_bridge_io_s0.address
		.mm_clock_crossing_bridge_io_s0_write                               (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_write),           //                                                             .write
		.mm_clock_crossing_bridge_io_s0_read                                (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_read),            //                                                             .read
		.mm_clock_crossing_bridge_io_s0_readdata                            (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_readdata),        //                                                             .readdata
		.mm_clock_crossing_bridge_io_s0_writedata                           (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_writedata),       //                                                             .writedata
		.mm_clock_crossing_bridge_io_s0_burstcount                          (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_burstcount),      //                                                             .burstcount
		.mm_clock_crossing_bridge_io_s0_byteenable                          (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_byteenable),      //                                                             .byteenable
		.mm_clock_crossing_bridge_io_s0_readdatavalid                       (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_readdatavalid),   //                                                             .readdatavalid
		.mm_clock_crossing_bridge_io_s0_waitrequest                         (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_waitrequest),     //                                                             .waitrequest
		.mm_clock_crossing_bridge_io_s0_debugaccess                         (mm_interconnect_0_mm_clock_crossing_bridge_io_s0_debugaccess),     //                                                             .debugaccess
		.nios2_gen2_debug_mem_slave_address                                 (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),             //                                   nios2_gen2_debug_mem_slave.address
		.nios2_gen2_debug_mem_slave_write                                   (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),               //                                                             .write
		.nios2_gen2_debug_mem_slave_read                                    (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),                //                                                             .read
		.nios2_gen2_debug_mem_slave_readdata                                (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),            //                                                             .readdata
		.nios2_gen2_debug_mem_slave_writedata                               (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),           //                                                             .writedata
		.nios2_gen2_debug_mem_slave_byteenable                              (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),          //                                                             .byteenable
		.nios2_gen2_debug_mem_slave_waitrequest                             (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest),         //                                                             .waitrequest
		.nios2_gen2_debug_mem_slave_debugaccess                             (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess),         //                                                             .debugaccess
		.onchip_memory2_s1_address                                          (mm_interconnect_0_onchip_memory2_s1_address),                      //                                            onchip_memory2_s1.address
		.onchip_memory2_s1_write                                            (mm_interconnect_0_onchip_memory2_s1_write),                        //                                                             .write
		.onchip_memory2_s1_readdata                                         (mm_interconnect_0_onchip_memory2_s1_readdata),                     //                                                             .readdata
		.onchip_memory2_s1_writedata                                        (mm_interconnect_0_onchip_memory2_s1_writedata),                    //                                                             .writedata
		.onchip_memory2_s1_byteenable                                       (mm_interconnect_0_onchip_memory2_s1_byteenable),                   //                                                             .byteenable
		.onchip_memory2_s1_chipselect                                       (mm_interconnect_0_onchip_memory2_s1_chipselect),                   //                                                             .chipselect
		.onchip_memory2_s1_clken                                            (mm_interconnect_0_onchip_memory2_s1_clken)                         //                                                             .clken
	);

	deca_qsys_mm_interconnect_1 mm_interconnect_1 (
		.altpll_sys_c1_clk                                                (altpll_sys_c1_clk),                                         //                                              altpll_sys_c1.clk
		.clk_50_clk_clk                                                   (clk_clk),                                                   //                                                 clk_50_clk.clk
		.mm_clock_crossing_bridge_io_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                        // mm_clock_crossing_bridge_io_m0_reset_reset_bridge_in_reset.reset
		.timer_reset_reset_bridge_in_reset_reset                          (rst_controller_reset_out_reset),                            //                          timer_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_io_m0_address                           (mm_clock_crossing_bridge_io_m0_address),                    //                             mm_clock_crossing_bridge_io_m0.address
		.mm_clock_crossing_bridge_io_m0_waitrequest                       (mm_clock_crossing_bridge_io_m0_waitrequest),                //                                                           .waitrequest
		.mm_clock_crossing_bridge_io_m0_burstcount                        (mm_clock_crossing_bridge_io_m0_burstcount),                 //                                                           .burstcount
		.mm_clock_crossing_bridge_io_m0_byteenable                        (mm_clock_crossing_bridge_io_m0_byteenable),                 //                                                           .byteenable
		.mm_clock_crossing_bridge_io_m0_read                              (mm_clock_crossing_bridge_io_m0_read),                       //                                                           .read
		.mm_clock_crossing_bridge_io_m0_readdata                          (mm_clock_crossing_bridge_io_m0_readdata),                   //                                                           .readdata
		.mm_clock_crossing_bridge_io_m0_readdatavalid                     (mm_clock_crossing_bridge_io_m0_readdatavalid),              //                                                           .readdatavalid
		.mm_clock_crossing_bridge_io_m0_write                             (mm_clock_crossing_bridge_io_m0_write),                      //                                                           .write
		.mm_clock_crossing_bridge_io_m0_writedata                         (mm_clock_crossing_bridge_io_m0_writedata),                  //                                                           .writedata
		.mm_clock_crossing_bridge_io_m0_debugaccess                       (mm_clock_crossing_bridge_io_m0_debugaccess),                //                                                           .debugaccess
		.ddr3_status_s1_address                                           (mm_interconnect_1_ddr3_status_s1_address),                  //                                             ddr3_status_s1.address
		.ddr3_status_s1_readdata                                          (mm_interconnect_1_ddr3_status_s1_readdata),                 //                                                           .readdata
		.jtag_uart_avalon_jtag_slave_address                              (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                                jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                                (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),       //                                                           .write
		.jtag_uart_avalon_jtag_slave_read                                 (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),        //                                                           .read
		.jtag_uart_avalon_jtag_slave_readdata                             (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                                                           .readdata
		.jtag_uart_avalon_jtag_slave_writedata                            (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                                                           .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                          (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                                                           .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                           (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  //                                                           .chipselect
		.key_s1_address                                                   (mm_interconnect_1_key_s1_address),                          //                                                     key_s1.address
		.key_s1_readdata                                                  (mm_interconnect_1_key_s1_readdata),                         //                                                           .readdata
		.sysid_qsys_control_slave_address                                 (mm_interconnect_1_sysid_qsys_control_slave_address),        //                                   sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                                (mm_interconnect_1_sysid_qsys_control_slave_readdata),       //                                                           .readdata
		.timer_s1_address                                                 (mm_interconnect_1_timer_s1_address),                        //                                                   timer_s1.address
		.timer_s1_write                                                   (mm_interconnect_1_timer_s1_write),                          //                                                           .write
		.timer_s1_readdata                                                (mm_interconnect_1_timer_s1_readdata),                       //                                                           .readdata
		.timer_s1_writedata                                               (mm_interconnect_1_timer_s1_writedata),                      //                                                           .writedata
		.timer_s1_chipselect                                              (mm_interconnect_1_timer_s1_chipselect)                      //                                                           .chipselect
	);

	deca_qsys_irq_mapper irq_mapper (
		.clk           (altpll_sys_c0_clk),                  //       clk.clk
		.reset         (rst_controller_004_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (nios2_gen2_irq_irq)                  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_sys_c0_clk),                  //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (altpll_sys_c1_clk),                  //       receiver_clk.clk
		.sender_clk     (altpll_sys_c0_clk),                  //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (altpll_sys_c1_clk),                  //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (mem_if_ddr3_emif_afi_half_clk_clk),  //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (altpll_sys_c0_clk),                      //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_003_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset),   // reset_in1.reset
		.clk            (altpll_sys_c0_clk),                      //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_004_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (mem_if_ddr3_emif_afi_clk_clk),       //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
