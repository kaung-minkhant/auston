��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��s������\�Ἡl-�y�f�����f� �ѕ:�nA�kb-q��_���ѹ(4�dê*���7��N2�ɐ��+ٞ�4Y6Mx�ejǴ�y9�����=���D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��\\�l�����r9s��@'�k~�{�<���y�#���i6`#Ɉh:^[����*`��Z��|���z���N?`q_���ר�Z���FLe���Et *�mkd��^�\D�{�Ѫ����+*����+�Z����� ��ԓ*n��an�7�?��!\�ݠͿ�L=,���a���Nk��_=���}�7�C�#T��<T���w�w��ƕ�_�m�����դ��*���	�4+��Ch�S� �-�6�똒��Om��9ד�0�XZ\,��zF?|���﬌62����&��)��*�GXW�f�72�!%��F�c�R[���f�s#U��"� ��b��*>zT�9D�'���l*j<�$Hm~��ˣV�=	ʥ�>�/%��¸"x2�hW��t��mK�M��-W��f��8������f��U"p['���]��Q����ќ���W#�U�5�5�S�
P��܁NNɅǶ�9���#�S�V���1U걒'zl�c���+���os�S���Er�����\:�'B7t&���ǌ�u��Fz�A>�J�rL��p�F�	*�s�C_�BM�僐b�Ĳ7x��P���QEd��d�Z���ou낕Z�i(��[keY�^��1}�".�������'5��+Ï�,�.�*It6�-��{�⵿��8?�C�FZ�fh+���oj������6����W���>��ك�L�"0�M[<���<��g��?/+��o �E�>��XY�ד�N框/k�y��((�N/%�o_�,��!���D1Č�����f�p�䔺�
���`#p��$�P)ש$�˿`��?k{u��/DP��_��X���0�&-qDǱ�(i_S9(M9��>dU+��&_gY�6������$H�)55��QK\�LD�$���cl����b}2�v@*��+r�����`�<�yz�����n!�9���;潠V�}v��7]3'�g�W��8�}��0�9,,$�$���s8L"r��qYj�sU�S�D^؀��d�;Kp���kUW��e�w3��b�q�o�h(��1���r�HP%1�%P�y �)�7.2��Yw|m�-+�(x�7/����"́�I��4�����}�>��k��15lu�&�1�,ͯ�-�OA�=]��"I��D��JK6pQ}��Ϟ���8��;�#�-��?���?]�����*�����L M&"�_���W��)c�����}~���!�eJ)=kN�����I�t�8Op�+>H��88ɂu(�����T�w�h+9Ah_�Cpm�M��˯�<� +�z��Y)hdNq�~�ΦO�j�z&9�C�`��+�0*����M�X-�������)+�� �@��M�$�CJ����OwIw4e$�3���o�#7ա5R��g�һG��C5�Tu��AIBޫ���;�4T����9Ӳ�
{��H�ڨ�;�>Q��A�Ҥ/D@"�����*�\Uɪ�|�<$��
y`��o��ִ ��w�
�����X4|U�
�^�p2�>n�6. Q'j���_7��ÑQ���=TC�·�zI�5\C�R@��b�N�h�������P)��$]$��TL*+E�]g
S�q�K6{2#\`5�ݷ�����̘]�9��L ����q�W�v�����_<$oo�"���H��/6Ѱ-/��O�u�0C`��M�ƅQ^���F�		�۳�t�*��\M���T�SA^I �T?ό�Y��"�z,�
t%��t�>�{��,�Ws9c�}�؀��Pj~����K��ⵯH��"�u:��;Y�>�S��\Sm�燢�3�A�C1���N�G��݊M�i0GQsx2�A���xM S�7r������~���| �O�����K�D6���d�W�ܗ
��c�J�f�T�a���2�céY�"bb^�3��R{���[G\Fۦ�v��7�ofY��q���+%|�[����zb�p��h�Vx�V��Vkښ�O�Pkv�;����P��q�c����]����2�	��U�W�]:��x���D�҇_�b��������{��������.�|���>��e��Z܈#K�[�H�2��@l�,���	���=�O���"ɋ{1ng�0@�6�h�6�0o-��o0��[*�* Z�V�䶇�Za}	C#d ۏa#��}����}�ʮT�Wϡ��m�Z2��ذ�"�B͖�tP� hx�$�o�X[P�@�'/���:y}/N�s��l�`���E����Rd�G�=�VbvjAW�md����Ts�L|�pM�׷�Ub��>MY�X�Ko�?T]0��\�f�7�8A��Ѯ���R
ו9>%��q��%��[z	$,�p��?���|=��wRPDN�TP5'b�O�'VuR�^�j��mg����o`Ù�п�c|��6DU�)��o�\Nd4Ǉ�T�)���-I�n�&?g)��1;S��S�Cx�F��7C���`��ы�v�R�Dsj>>Z��J�8,#k�~K@2��+S��GS4�%���G�vC�nx�^5��D�_�F�Y[��F�r@��#��,�e,Du8���(&8
�Fu���P�`ȯ���m�0�Ot�Ļ����7��J�&����h�h���8�u��;fe2d����°�s2x��r6-����$�v�yB떚
���.�;y�}}1�ۢ������ Ԋ�R:�R��Hշq�'�Q�Ҩ,q�UG��,PG�:�V������?0�_k��f��2gن�i�͒$�~�A���MGz�R�8��1�uꚈ��gL~�}��a�(DhD���.G�s&M��
FԍpD6�ẹIz�,+'�(�uΒiej���Ra�8(�:�9����E�ӮA�<N.�	�_8�{�2�ZTP�G�U��s���<�&ER�y���%�5����f}K�s�ʕ��yn�{5���Ж�V�W�葯��8����*�Yƥ��,
�ご;��2y��i��&t���u_\y	�F�o5&(���e�q �0Y�1=^	�X��+���?��,���e_T;�C��; ^�J�&ނ��}R�	��/�q���D=�1����zh˥�C����%��E? W��s�P?��-�M�����x���hs�:�����<a����C�VDFmS�O��1RJSk!=�)��N�b<T?�	��|�vϯyI��qz�	�;�ױ?�O�����AKK�H�+��.�VvN~�D&3� VAUW���b'{̭���b-�&1,��]�"]��Ў���D'ۂ��E��R���^��9���5�ѧ�F)�A|8��������j���<�o[@�y/\��)ꖠ���r�%l��fKTh �Z9`�ps�K7��%<Px1��^�줪�j:�4�1�����R4�qݾ��iQ7�k��
k͔y]���ӏW9V����0ih�[�Z�U�Z�2���H��JطG�����|/�
�L��!�i����#�U��=n[m����C�Q�G���&�����E�f��m�GOs��|��fȤ>Mz[]�0H���-�"���A��qA�2���=Tq��,��V�i���V�ل4�������Pu�S��<�f��^t�����Ց������� ��9��eӲ	�k纲���v�[��3�(��~�����l>��7�P[���˖i~�OW�~�,�ƣ��/2��l]?�{��G{���q�w��h-�KT~��sv��	
YG�-�W Ų0ص��CR��R5��|/\J���3k����p��k�Ӂ�b��"e�I��r�*�h�'�A0��ThI'gk�8��ڽ�|	�!���M����0���/�h��7H�֜�P�۫Ჳn�����z�J�0��NE|���8M͑�������u�Q�1��s�4�/U9JY~K
p�N��<����om�����]^�������1ȕ�Ae�B]��.4�ޣ-��%Y�@�r����[LX	Z�"p%�/SN?���ƣ��g/�m�����bݿ�e5p���j��Tߛ�Ѥ���YFi0!H�	����Ygp�%�(-� ?��pM+1̝I��#|G$x
����F�)k�M{�+��T0��K�ð���{a�.,����q��S���MM���S��/�0*��42S�+֭Vd�l�31+�V�kfu�2�1�lf�K[�IE��*}z�IjZ�"��oxo�gx��~J�ꭇp6?e��>���C <3�VE�4�Û􆳷�l5�I����kt��a8�>���Vïz�������&��_�Mm@ˍ��|�T�;�̮˞~�2��ʢGղ`�`хG"e� �X�Nv$:�c)�v=�p�݄����?O����ۆ�B[)�{FO�U����k%˯)`��sԓ�r=I��t&$��X����S_�U��;�zhģJ}�V�U�Ť���a.%�$����}����}�W�v����-n
SZb^}�q�iKyAi�P�+,ê�[T�엩c�|�wI�`�''�F�]�MޠTY���J�vF��1�MY�d�*	)4��zS�+���|1�m~��L�aqBo��;��p��>ͷ�}#���'v�o MB�[���w��%;<��_RT�}�[��F��r:GA�
��i��of����er&9D�V������i���ԳD�:�����$�MOۮ�k4�wV�c�}A��*�i̫CS�"�[�͗��y��M�����%8���}x!h���S����w5���SY5��<|��n�?�Z�'6En}��>�4���1ʴ�ya�Tf#��� ��E<:凉z`(�j\�ׁ�C��_'��/f�{H����8�q���P�bn�$�_I9�ҎL����-���]��]添U-*�FW�@`F�H���)�@��{����u�+쾭��t��u�cTH�}���f����ke��냛�)�QM\��F��Kð��/�X`+FJ�����ܮ�%��H�
�t Z�Tjaֶ�������(��]C��ZϢlp��FL#J�w1�:00K*�G	�ߺ�3O���3x������{��$��g`�A���m��O�,��4�A󹓄ˢ+'��oF�d&Gߐ�sC�0V���+P�"_c�����жi_-�H1�i~%zƴ�Py���FAC֏�	\�/��ԓ����/�v����$T9�Q���$Ĉ�-	`Fh�U�Z���e�M��o[C�?�:gU��B�z�ֹ�P&���;�5��ғt�,��	��^A�s�/%�P�_�H&KD2c���$�ʸq��7)��FNMi֒c�E�GM���-��%O���֐1�Z�Y׃(�`<�S0�w'�b��e��E��ϓv�4C�����/О2��~��)v>B0*?Ġ÷�E�[�U���'�<�/�-j9Q�Ϡs��M(�<G�C����)��bx��wA@hHE�h�l��]H��]#�ۋ ���\]S}�>�z
a�S4��-Z;>_��h�����z�P�2��/���ÀX��2�-��>t�0q|2��p����Ji���_so3�Fn��V��`��/�O$�<L��ٲ-���z�ܧ8�8�JW�>=5�g//�~�>�ΣIX=^F(�ᵰhe���60�B�<�4+��t0O*��E���d㙮H�����	�2�j���8�l�UkI�������D�FF���������(CK�a���g5j�_6��w��۳��^�(O�GXPm��3�,�M�3�yǥ���j��Ά����k���m5o��?<e�{B�U�)!Q�����8�c�o����SKt!A�W��^���~�*��o2
��6�` �~ �$!E<�+hږ
�q}u4D᫡(���Y��bQ^��q��к�n�e�;I'���<$%�4������̳S�c�*�#q���v��� �_}\�
(�O*s�&?&��]����glΩND�W�W����!���c��r3<	y]����\D,-�1�Q��;.|�Tv�¿�&@����U��� ,��~f����]ZQ�`����@� �M�{�=2(Q){�ZBcg Ύ�JLw�y���yYU2t6�����A/�j�f��]$^N�?$/���kfU��t��_����xeK���۞D{F� ���Ɗ(��D#�0]�U�æ%ʏ�x	��~��N�كR��������a� i�$}�R����n��#����J��m����򞃢���N���qc;�?K��N4_����L���pl�&�섙������:=3ʜԦة��#�w��j�����A��,	����s�2�tO���0F wp���s|����F���=UM�l�aX��Jp]b���������Pc�O=	> IRa��_�v��9 A�O�C9D�ee<�V��\��߸4�/�����m�Æ��)����O���	q|��~vPm���v�@.�=;ga�4�>�"����q3�����R�W6ٹ�y���F_�/]�Z�]�co�z���ZΖ�T�z��i���W�R�S��/_�(����D4�������B��g��z�@E$�${��N���{�+�(�в ��m��a���T�r.b��O��i�@z�}�W	=~Ӓ��4"��Bʝ��N~�	�?$�)>�fH~�!J�U��T�Dm���|vZO�̀~	zː'��<���ݑF�����s���)Ք`8|���Q( ~�qu�6ƭ/��U%F�}����g���j��=Z�k����U����ߣ�&cY�2#T�1��y���t�+�܈n�4�ۄ�J�1�iq�.Q%�s�L�݅��_�<?H`��?%�I�p2��2�_M{T��BΨ��a�g]+�����VQZ(|0����E����H3
���٨�;g0g����nK�����?��bSlr��]���l�q9h���Δ�=���	�2Zt:�Y��$ݽ$�+]�P�!��b!�u���=����huW�N��͝���Ʉ������&��BM2L��jh�Yg�Y)[���/�ɻ��=&s�����GP����c_k��?r�t_�%@d6��e�~ۇ3�?�'A�	��䃛pa�������fX�S�X[��p5�@����B��t09ť�a�6&�Y���X�$.V}�#A�<��=+IrL�ԙ�Ѷ����.�g���!�S�Eݝ� �t�3���w9���j��]�8��7ps޳hn�}�kEb�s~RU�ڜ+�K���l�S��K�T� ^	}3����uq�'7�T5	SW&*T�L\�\)��G�P�3|��b#7d���n><�����������Aq�>�*���F����ٟ���c�P���׉�����*%c؎.s�u�F	�פ�$д&��8���y�6�k`����@Y�/��4��8��
̻�P��O�����a�*�w�=(��D����ǹ���/G����������K@4"�9��ͥ4%�	E�N�h:򍨊��H�̞a��޻����.z}�_����Ov�8ā�$d���+�����Ǣ0K� [����8��/�<T��*MOp�]0"�19nۘ�%�U�s�}�0���w_Q}ήm�ǌl�i��k�<���<��>�!��/�˲����+�Q����(^�$�R¡u��>�({	��^�>�)�����(^y��*�#�U�@LKQs��5Aw�24W����l��{P�z��k�%�&≠(����V�1���h�$��Y�\��]�&��DŽ<��3�~O�05-�:��P}3�A�s�*�3�/Ư����E��� Qgs��ٷ�b��o��	�K�� ^��Տ��L��	ӱ0ÆĴ�U����KQ뢎���8��������MT_��T��/�B�{Ā�+���u�4F���(�B��'���pcÍy��=�G�I�	iuȢ��[��G������6
宑b�idQ��8�յ����x/��?Y��'۳��UX�l8��4�`G��X� �0ܩ��>��~�M�����mK���>H���zȭ�@t�]��]��e��>Eޣ&��8X�9٠��������� V�x��F��L��pl�N�FW���}4��� �4@B��Nj�IUD���y=I�%����J���;{�g�zkO�Q��x	Z�<��
Y����7��Fr��*bp�!�Z�^�%�b����̅נ<�ߔ<ei�6��!!(\"W�׈�n�ݙ7ͷ̮)S�n����DI�"^�G��BR��̧`���hX�'��ٵ����jwWj�[��ۑ���Ϩ0�<�:+�~�b���Z��/�^
�p7���'Mu�=Q�wzM�g�$$()���?�
�AM�,h�PEmʎ��r��) jI��u&�
m���1�������e�_=�`k�p0�w�Q���%-��?���1s*ܛ��� M> �{M��j�^Z���E��^�2��v��1<���I��MB���1��RT`��E����a2���m;W�4n��n���c�&,�R�H�P͛�)�1x�;��0Y������j��d�[(I����R���u2W�A�ٰ������I���n���#�l�;����q)z�`�
�N��YLZ���KJ�����M�U���3�|� e�#�����}	�J�6��q>���C>�Ӷ��Z^}��k?�i�S�}�4_��v���q^:쟆t@K�g���R�L��Q����gr�I砌�κh��Lev�)�����Nk��;�8p�M^RN� �n��x�:͹}|�Ԟ�z��������Ĩ�SMC���7A
��Z�����{��_X��U�2��|��P�t9�܊��S��C�����f:�o�~;��"Δ\���s���(E<�,pi h-q#h�y��?^Bֆ�~nnJqM9�:<O�6󆬦63t�1N�fTC����F��	���!yP�R��T�[<�,K���d(s�qG.U��c��%�n/9�駉�\9Tkm�B�8徃���1�)0�W��{�g��5I�L��^�հd"ڠ��c6XfIXT��r�'����BX@з0�+�߯^Ց�a��+�+_F�mF;��J,��0�H�0��3���]`�)����T��9��^���$(a���T(���f�Yٓ���{zІER�m,�vL\|1������?pw���uO�[�߸��DG]�}!Y�
'#�f�{���F��y�l��@�]Q�������Y�%�����5/��v���J�g?�$O�P�js`]��	�ݣ�N^d��l[Ćs��i���	����r���8(���T/��~����|o����[�
����1R%�d�v��N���Xu��L0
������~��\��p�������[b����[_��eapu�y��R�=tV�!L7�T�����j�!AioLG�a8ɯ3��W����魜��#XAyix�~	U�""Ie׵O��f<Sl%֢H�3�}�NW\�*�ڪ]�#S���qfin_?̓Z�{k���o�_��P���`�'�k�+8,kw?��:bE�*
��A��V��!��,�d]f����@��~y	���E�q��j��;��fI}\>%���F�Ã��+=_�z���W�s(���DW�w�V)�j^@Z+�D�[O��o�sI& ���+%p��Zlm]HҜ9��,  | s�{D���m��M��Y�� #��������`�Ù�Rܕg}��>��9ź���!č�`뱰l
ʮ����4G��Y�Ntb�k�O9#�&�5m����*�>ݰ�E��aRό���uA'�m�Qr%�C��Y�Oq�.J�������
�\S,Ɋ��m߻퐸��E��Mm��T���]�ZQLx�1��@�ZJ�ZN��s��YS��W+%?��>�niU�9�������):�������e�܌)�+��Q�<yt8���ڰ���É�H�Y6�3^DC�/a�^�$ܤ%�0�lx�${NBv�p���Bh1�f�++V~��r*��'^���u�����f����j�̊��WT���ݒleK�Z$���R�Q&��}Ky��2���!JI�l�%&��p�ۇ����;Kqy�!��^{���?oCf3��'b��Uk`�e��mE}WlJ��9"�o��N��&5ĜȌ-�~�;V15���� �ӧ`$�IW�&��fc����m͊�,U�Q�\���G|��M�	:Rh���Mèi�s��/�-�_4�N�T��x
�m�c�RqxJ�$���w�!�F�P:K�r0YZ�:�m�Y���{��H�����&����|��{a��OeF/�-���p����r�k`��.V�YlL��ݷ�BY����AӅ����_�u�XY�8���5V�2��x��W6�Σ_@�c o�~�T�λ�SlS����G��c�.��O���6�{�ܨ��Q�9��|l��:�)jVm���'�D��!�q�d>G/'vw�\$��F��
������֛��%.[|J���99{F�Em�-0p޾�w�\Q0ڦd���8�aS��ӣ-�Ȯ�g���v��
m��ݼ��\u��H�ƫVDN70��D��ޞA��21���j��o�}�/�ZH7<ʊ&�+"P�59���J
"����#�E]�W ��Xǐ��ַ>�T�0t}/�ě�	�@O�SD�Vo+�_=�F%��٢�b� n�s!@!n-�٢!�U��<J�� ��ӴqMwj�$Pe(On�$�x�#����P;���;���+��(g H�]���ֳ�Me�3_Kh���b⃳�!�}���-�l�ϙ�(��:((��=�%5�ڻ檞��A̡}���g��>���*��<��RJ�xy��8��ۥ��i+��^�Z�ü�B�+�j�D��5|�����K�Agt\.��3&V�sw�,x��u������P��I�oz�0ٳ�{����n�I|��gS�X �X�HN|�X`$�ȃ[R<�G��.O�ȏ兔b+��C�g��5���h�0h��\o�<U	��ڀA���9\����3�uoa8�;�@��������ais�]�rc/�^�-���I��Aj��EU�%'���dH�,9���
�i�4��� �>6�d���J[Y>���#�ED�Dˣ'������]z�d����A�H��W�sUJbV/�����V�M�CU+�/,t8qA[��n�P�b�GM�zEB�ň�^�:T�T��=�&_~2��tm��>%υ�j�کc;!��ؙ�����șN���Mh����D�V������C��Y)>���Ea����'E�s��� 7�\(ƿb��-�P���w��ϖ�(J��[#_I�o�ŜY5�wO�`uo�%�2�d�N�ͬ�yH�vC��8�Tˠ�?
�zu��h��F׺\�#
�-�c�u�`�9�L���FI*>*����ˇ���:Q�M)E�34[Ҡ�Ix�58�N'��7p���8\\��qx32����<���b��WEG%�?R_Қ��]��ǁ=����5��w	zۉR�𥅼ǣ�N�n��HhF�)ϝ�*�燊�~��K�nB��%�g�{�T�K> o)U��xV&�Gt�����.j�P�K��L�o��n�P��w!�wze,�}%���+&o�[m�>�!�<y1r�Z���>\v#ןzQ �XP��s��x�3��s<,��9F��]��&��c�=�w�iG�s8&��ݍ:BT�k�]��m�U |�)5�Ӑ �7��[Ԑ�W5�Ǹ/>�lC�Q赝�?�9��=�ɡóG�j��`����@s�i�Wǽ'�خ�(U����v�ێ1�^:}�Z�r��V�^�E��ji�����E�,`@�z�0�\�h�5�|)�ױ&�Ab[��鸬�����-I�܃4fA��?>*�]��X���j��VN�q�6j�^3�!~��o4A�����[�D����ez}!��@R�~"n!�<�0у��O�Zh~e
89�w8�2Hf��z*S}�����c�p����d��;�y���0��@�s ���|zU�6^�s0�,�$]!�6���T��X��X6
7���U&�cg�+�HC��v�����s 1��l#�!�3�+�|�)ǫ�vv\���v��VkS⨇?mG��$`��.D�z;n�����@��� �ą?�1�q�*�̚��8{�-�CU��Ɓr���{!� t�Z�ێ1�.xD~2�jy}�nO�2��y�N��/AS1���x�g����`h�4�i�k,����Uڝ��7������v���Z���.0i����{ޓ6Z���Ҫ��XH��|U��q����w]1��QG�F��O�B��{[�>t�"���l����n?��nw��k�߼Q����Ԝ�̈E_c�CU�ݾ��^�#5H�<A;l���گ�H�1�K'�w	��^�>�
ͣ�;S:i�n�Ր��*uG��%P�	4����f���m)�҄C���M-n@�o�Ӥ9�.)�y�#��+͚�����a����!�k���o���S��;�l���l���Q�Ѫ]�f=Uk_G��Z��If#y��m��އ��ST�.����D���oFx���p̋�����7n]��GfK�&y��\2qe����텁�@܎[���'�� �����=F>��T�[C��{h�2���&��|b�;�x%��������	`�Ɣ�V<�����=���}��"�X��;�Y�e���f"?����}@�gJ�\J{X�bUH��k�'�b���ͭ��g�
��2�0��Q�-T9�*�o�d�Z�Ĺ"
 �}�˺N�& g����U�R@j;��W�F@���(�{D��	e�ߍ�LPE�~��1���w���ܬ��T�A��T�,Lq2����$�˫eg������_B����m�`��3�u69��-y�ƬI�����O0Չ�p�[���q�ل�~՝��:�[�1=��PT7�&����7��\D�0�w�;��i�F��D(Z�)*�U�X �����!9bj2�O�{�ъ���el�1+3�ٛ;^�
r/Oo�՝�\�zS_�|�W��I1<�;%��،hc��B��d��q^V���Cx�S����@i��rȚ�6 u���F�?�z�ES���j@\YWH���#@� ��]��+8z�l����Upo�Y�H{�`	�f|�:�*�<�E4������54s)�Չq�G#��nyb�ts�zk�u�Ƽ`թ��=>���5�Ģ�k�p��P�P�2�4��� g����
o�[c"[q��|��C;-F�yΩ�~R�A���_��r���ܔ����D��3B�~���'=���3�f5~���c�T9��W�23�6�V=M��FZB�1@Yi}�N�~��h�M:2�I��P$�z����SX�(��qW�[1Q�wޭ7��_Q�Js��"σ�i��co�K���z���Q���:�5�o��c>d��x�C��:�wb(���l��}!��ц<l��0��_Vx=kP���ޭ���|�������,�S���z�ҽʋ��'���W��'�:�:y��G�P�g��~�*��&��-�A���[� <�̛��ɽϘ{0���kHl"��&3��_՞geb�Ý�Ѵ'��#<ڪ�`�?oT45h,.�Ӿȍ�y��m��G��5�OYɴ�O�_A����J �� �b���h���6��T���"�I_��G�:�T>�(�x���%����g/AH�TX�U��1��P7��WRV�,�q��6mk&*@0:�1H�6T,�WƆ���<��8J֞NÔ����%��O���6c�fI��M��xU1��(����[4�K�6.�4~�TA����VR/�,=$�2�XP� �.�P��XJ];���&&:�ݳ�����!?}��De�����Υ��Jr6<�an?{`s`4���{���E^�
����Y.�V�|���<g��Bݸ���e�*�ݩ_�$�+�MA���P�u���~���IU�Zp�r�)]�>�w	�`�h�/�r���D,Z޹?rF~���*��y�;վ��	�qS8*������Έ$����Xʕ�Ǔ`\�^�o�7i��4$���L}�=��^� ��$�wp��NԖB�[��Lٛ�t���䈌���'_���+b�H�F2$P	����;¿��ϒJ ��;3j�wY݁O���P2���d���Tc,��A�C�NZ2�A�������Zc$���h�~��5�c�]����Ό�$�A�N(�:\��q�q�����77���:����sq(�M������F�k��.&Ƭ /	�������W%�>��R=��XQA+���%)�R��g=<f1�y~g�M���1yE^zD�=T��谬�ͬ�s�o"Z|�!�W�Nj���5Ig��M��]�_��
	��N8���m�TC��GT�<�@.T�&�W�'����H>7�L�hX	�tMf8	�)n�S�V�	�p�<��AZ�~^ԇԁ�˹M��%�ǌ���]��+��4��F1r��v�K�Ht�,K�.�I<��s'�u��O��� O���ʢG�d,���T69��1�y?�f����kQ����G���1֑R$J��u�(��H�.V9��E_̎�F�؞|���tC�`z�)v�R�FlEh��{H�Q��'���K����kDB>��|�壣m������W�IO2�֤�'�F��}�)���Cc<r�l.9�������+=!~���|[b�#j���db�"���j׈�J��Z�k��0)�Y�ۥ���ְ�����6��g�5c7�z�v�޷ U.(7l�%`Y������(~[���Cj��27����g�F]��CL�&��H�.dv�zXu��۷�^��Wa�� �F3˩�*@k�%�n"|
tD�[��:{W�^o)��9f�������j.	e!"��Z�.��}��N����{ץB�'�I��_l t@��ĝq��/R
��Ys�cҕ�s��7蔐ˣ���QMv`�qe��V�<��������}��ͷl{�'â&��ۼ��M�j7�nB��,�=e��d��)���é�)R�b�v�ނ��'<ч�P��`��@�X���ګAȪ˄��$7h&:jQ�p����E�����.�����<K�Í�i[+F���g�F��H��(�ŝ�≽V(�r��#��`�zh?��h	�0�gGO��F���d���./�bX�(5�?���K(X��Ws�ۀ>2� �H~�Ѽ�?��+����Č3P~� +�Wl�ؖg�y�R?�^ё�R'b3��а0�Ԅ�@$� ��3;���kN�{!�?���V��ĵ�;}�;���c=}I�����Q}�����+�-��CE����5_<�f!-�C�M+���R�
����*WGty���Ҟ��8��� ?y��q��u��>j,(��; fm�\�j��uF��'Ud��L(/md��)�NٗXF�H�x�
O���^3���T����){.L��A�� 
�"|���-Ѳ���A�v��,6P���3��4%���V����n���	�^�Ns����_��H�6�F@�2��-m$2���Ljڭ�]q*�� c���\K��I�u�K�i[�����qk������<��t믍�ÅI��WgY����DXm��r!��g��ܵj��\��0�\b�����7>tn6�AG.��l���O�req�K�>��p��tֶv[�s�(�.��u�(�z��ԕf�.�|��t1x�]��^+^˃CН{�q�\O@�еC�F�1���^g�J������C�2c �R|�P�,w2>���%��5߈���;������p�~s��|ۄ�Rb:Z�Q�_U}�בd)�t"áTY�b(��_�R*'T+߆����Ӆ��_���ث��\�E~�n���<��`m��.pS�< =��8!����w�*�]�G�䳌���R��h�`�/��iB�.���J��a	�;�{wc������O��\�/"Xt&2�B���ɲH���6����K�?z���mVN�`�����w�]\]nI�Զ�ʅ6��Xߝ@|E)?�fnT���M���������=��z�lޱ�ڥ���=	�nH��q1��b2i�3���X���Ij�%P�%��ݘ�x�{�D���DA䮶0���y�4��;��!
M��L꾀�x�+8�Xx����aP���$ގ��j^�Sv�-�O|�w
ֺtw]pI� ĺs^v��{'��is�nE-�> u��ܲ+�.��Y���(f$O3G>$�������K4z��;Hd}H��=��WDM�{�����D����N�H@&���zt*�|g�%� �N���#v��zI�.j����,�A�{�zJ����G��M����s��W%G�� � ^Q�TYȊ%��)�[ �^R\;��%	�pP�KW@���k�����zH�\
�����q;O���凒�Yl�#����◴���f�<^.� �kK�J0�� �zO-�#u6L��,���iU�_��ħ|��Ą
ɆQ��fPr��Kr�NR������ �����$G�NTݮn�Z0�+/��oj����� s���D�w*�zn1�������3%�"J��B
�M��F"�F� ֿ;X ��	bO&73D��/�;�=:P��V#��Y߮���2�]6|a4���Nl=@��A�ț���b�Vh����sol�:�X�LDx��z���r��K�?^��h}D~�eHL��L��ƄQ�"��se�Z�-B^�_�`҇]���S��O�6�zz((���Ԟ�C��3�^���"tB�.������pw���&�/�\u˭V�5���(�C�mjMv���7j������z�����> �.��;�Q�pzf# !�*j��7�n��@��\N�������B��|��ա�p.&U����(!�Z��¤Z@�?I8��
_�g��!Rl�햋�H+�J�@��؊"]��v$�ΧI�{���$N>�~�Q�q�^��G*��L�
:'����e껰[���l��|��Wd ��$���k���ՠ�Ȓ�����dQ�3���>:�4��xz��`�����%�����_���.�[I�!�W�_Y�]�6�	�7��`L/��\���o��T���8�h�O˪���|ǝ��{�� ��JqI͌) �d�]���4y��ȵ"_�'��O���	�$"Ja�G��0���d1��_�� &a\z�6�:�6���=�'26{Ȣo?�7n~;�e��H=�� d�(��dI�]���3��1��`��U�� �)�"��Ul��
3���Q� ��w��啴�]̀`�s\�IU�(f�[M��x���D�)aXE5B��*]om��R��-z����z��eT�Fm�2��nc� ��m.G�����x>�_��;d��F��>[uV"��UϘ�f��/����c���]d�{H�`�h��S�j��n{��J'�)k��`:�{b�6�^J���Y`N��	s��Dt�Ww���Z^X'��M�T�͠�V/�(.K[pk�b����
s�-s��x����x��h��8ti��}�Zbt�/MrS� �9�(m�"R�R���@(#:�?&�g��O�� w��g�"�b�x���s�/A��^�l���N�FAB4�ܔw�u���_{�y6���m/�0s���t�;�� ��KM�F+)��4�������0�U�Zp�"�Ҽ�{�{h��a� �����7�$�yG�ↁ��K�_��zk���Q\�B��E	�7������>r�N[�V�|`����``�!+\�8��W�ϻ34=ظ������K��L�Ҿ�P��K���\I^{���u����]�w抚!�ѳD;�`{i ��Ʋ=QΫ�ǲ��Õ������[m}{�ulzOa�����ȣ��]Yyܫ�7�x�X5�>" �_�XzV������=�"bE"n�Ƶ��:�<j�Y�lCw���I��1��ZE�%�e��-�zܻ ���y����~��!�d/MT�i|�8����YA�Cf�a��g��u8;:+Y�HCZ���y�p*V}�9�}����,�P�B�;]Z67�
���gj��w�8�w�>ck�e�l�La�dOB|У�zT��h��$��Y�渮�&v$���z�
����##<Gq4��FG��$)��5K�~a�n}bƢD��)�+ж�Ԧ�Ҟu:�[mp��v�F�E �#X�d��	�K��)_�7
NI$ҫ���w����R�e���!����4������Ꮓ�:F�]s7�qBy������:s�j7�w��3n"�eLMb�v�� ]��y���2΀���}�J�p����x�u r��*�س�J	�[��B)�_Kw�ec����r#��5G�����[^?'����W�nZ������w�F/��� N�+��U|� '!�������'��H�"��z��[�J�����_h#_`�, �XZ�����K�I�V��}4[�o�~���LM�q몮��y�,���^�m� �O���`  �UNM��w�_�p&���{�YV"ݸS֗�ı�x�û�������K��+w��d�P��-�Z����\�|b�x ����b2-`�oҪ��bKA�g�Vi�n]�6�����4�%+�vG�F�v�	�*���z�#�`��qa��turz��˖�ih��o�?��\�i���m�ck��	$0�?��s�^�d'��/�Y�&��}�P'�e`�z���X��v+����6��w���r}�yaxP���jKܵ��Si�`�!=D�j�&z�+J�7�MMc��L{�O|;;�>Y5Y�j���q�0e,� b�L�O�K�+H��J�g&94�v}e�L�"J�#w����e
��> k{���s��֋��vx5�)iWn�B��Zm�2�❿Uԋ)����y��7����& �)��+l
���Y8��O
�#�nf[#�]�ƶ_��j^.o�ǔ���߇�|�����h�Z���]&[u�Sd��y5����E`� S�9>��h��5X����64��+�,�m.>x"�2ѡ��w�����J�q����뙑�z�K���a:�[�m�ɿ| ��+=<<a$_(��LU��>�P U��x�v������!�	&�Wl�j{4w�Q�������\(�$���0�Ι)��jU#�/0�~��^�|�9��#Eks�$�rU��|j�K��N��V��ln�͎:��TU��۞&.�: 8<`[��$�����.q�����u��%20l�Lm+m>s�JF��v�_Ӿ��x3�	�~�fY��k�Jc�1_6��0�f���-�B�|+�����;��#�&���d �o�-����o���d�>Q+B�� F5'��aQ�K�ъ�`��T��Q˃4Ҕ�h�
N�|9�* ���Zs]4�3�p���6��<Q^a¬�O���[�E(`�!��K!c��D+��F[ث¶K�F&/3BĄ�#�S��p�)�뻧p�/�޷	�����M�H�������R���i�a��u���}���c��w�?z�[Ӯ�~Mpa��Tn��|�Z�N�� �?Ln������N��d���M^;��'��)�a�k���*���Yh�y�v�j�+1�C*M@������r�!~4n3�hr?�pK�V�6�y����0$s1:�=��&U�v��z#q�B𡘗[��,q��y܊e��c6���s?��4�^Wb�z���f}M��K�&|��I�`�c������F:@1����d_��|�b����x���`���)c�7��1��P`H74XȬ�hMx"CxVX�BL�]��!�#}VW�Dù���� iIS�$���X
2�v��"��@���@�'�'�XCfy���}	?54��(5]����[$�8�;�zu�%�����p��c�qˬq[ғ���$)�5`�{ד��VX�︰h���p��`T(�L}5�¦8����˟�V��[.Kf�M���CͩH��ȶi�(oy�r�x���k4{�JtJ�a�J��L�Ի$YT�v��n�[b��eQ.�ْ���b�������U�!sz��`�
�vن�Ȋ��m(d��yˇ�� ;����.��!��</P�:t��1j�煞��ɍ���m �L�4�����}reH <�J[-��9����AA�^~�����;zޭ�r뎌JMYzH!1�9p�d+��9U��h1r���o�]��8/d+Aج��0>�����)�b�2)Uh�3�F⿁(f�@P�d9U�k3����i�00o��C���3��]i� �uTZvN��*�-`Q� �����m� p/ͫMmv�G�Y�{�9��&�Ȁ�>��#�E\XH˸�����E�I�6j�?m������51����b�u�KU��g	/_u^YF�"M�Vo���Q\Z���\�����&���P8��G����l�M\\]�R���'�8���J�����G�����' ��(�}��Qώ�6T!3}��~����EP�}����iRy���;T��9��̿��/����7'������5�_���:_��`�M?�W�DK�Ő�KA]Ѣ,K��ڨi9�� �H�?zKv�5z?)nuZf+�o��T�I��ohO�Rn��H���kX��āH��e���Ⳡ ɳ���D�̔}���A_��[u��p� �Y�ڇ��X�3Z�K��&�OԐ�A9��w�b�,)�VUa�m-5��P��ݧ:�2w$��t!�i��=���x'��t�.kB���!`�1O\\b<�+�k�{�6Do������r]:3w�Q�/	�,�I����j�	��_I�OԩA�C�7'��?vSuX�䣍%˥&�d�{�y-�u-���+����-�+�-+َ
������rX���b�y�qa�;T.R�Wh���Z��^�����U�o��b+[4��w�'�?��p����x���g|��zl!����.6"gV9�fy��/ΈՄ>Oͳ_�J�"��O玚*N5�i��8b⚔ �B�Yd��yi��vǊ�c�X�RJ�x2˙�|M�x�ѷ}6H�������]�}4'dպ�����;$�}�*���3���~vh� l����O�A���6�;�uM$���>2�P�pn2U�$�h��ؚ� 5`[߷)��TpDp���_��b�\ߪ�(�3����-����P�9�����?מhL�v_�\�㎫��~���C!o#�f���CQǧ悈2ߚ�Ż;2nJ��[S�r�� �n��a������0: �M%D�������;����}O@q������h=���`6������'`g6o*6�HL�
Φ�b!�(�ї��ױ{���t�&�I�m�@d����9@��1�4LT5���o���ķQ�7E��{zף&X�PO�;Y���?*�Id�I���� �2»ڜ�9t�kMpb.���*cG�˨&���eeu �,�j1��F������͈���g+�������E�_)�握���p�"[N{-���36���/Kf�2�x��P4(]��l��]?�Q^H۴��{Z�f��S���Lo2 t&1���tY�0�!�Y���߰�٨�6�JL�m�>�OjA�PKh���+��Rl)=,�v�n-3`�Br��o�r���&0�$����M$�5:��Bf�E����/;'/��N9�5�X����6��'�@>�?_�z3/-����Ĥ�VC@�?Tֵ-��:q@��v���kl���+�[�&���f�S���i�2�c�إ
��n4� �xyÀ���	�\Q�[?�Pܼ3�bN'N��*�є�j������.��Bp{����`��)�ܨ]�}:گ�k�&�F�F�U�4κP��(?�-2^;�/�5sk��=_~�4=z5�g�o���A'�
B?i�V�/�0�Ql{lEr��F�#i��!�Zoi�
3V�����'%>�P�BnVbJ�#�H���E�� ��g�����g���a4��i��Z�ʾ�2��1�Gr���N�F2?y��`�̣R��� �{�!�gK�Q씞�m`b_�q��( 
�Haj	a[~��0��Єf�\����Nc��djJ�^Q��v�D@��qY����֙��۩Y�cV|r6k���̋������,_����f�UU�ay���îT����Ō^B�AK�}�P��C7
딶���>���fA拃!,�L��F�J�4��-��j��ql�E^țfv�p�m�݅I���<N�v]"z����U��'���u�J_�HZg�6ik�-07��s�����=9yށ��P;�����tﰻ$"���:cy�J���%�j��>�����c;W�$Q]�T�� ���+t�O�����~�8��L�{����x�A�����Y�1���!Z?���v7��ft(��}���if��Ӻ��x\!�
�¸D��@q�B��&�'(Ŭ]�Ms��[;���+�C���N=(D�M�!�Я�1�;��Y��nb�oQ��]np*��E�@��Q��a��8��6��-�CW��1����U�/���q���!��o/&��͜��]'���,ǒ������ޢ#R���w_N7N�=��el"�ͼ@s�Q������;;�	Y?��B�-�v�('6����Kg��Ɯ��;���Y��a�:9��I��f�^}�F�h����
p�~�E�!}&��q+����<�p8���ܝb��4�
�n^��Ol���=g�G6n�s���i�KR�@p�]�
�\#�39��~$
��ix��1��Q{�7c�R��2v�1C�n|� ��eZ��9�� �KG(�D��tT�`ڬ��e��Q��F@�E�S�A�,87K2��mɝ�Rd��vN��u�$ŵ׸colI�L����t�m�� ~M&
rŝ�����M��/<��P����d"���=ХY�Ģ���x":U-on"�6=7gc#�8 ��
��k����J�;.l:�ܦF��'�33�r�x4��x��,��T;$�J��g܋?��$�ڕ���d�$�O:���~m�F��_,=���$����}�H��S���NQ�[2���h�r�/p�`He�0ļ�����/%N����	�kal˧MU@����e���+���@J7�� �>n�)�nk�y��
��!]�u��X��?�w�|����FS�#,���E�U޹H#�SP�l{�*����w��>�B���N��o�Ҝ�̘k%�Rt#�=%��L��Un�m�U��_�1�v�Dc�$����e-5��1m�ưN�<��s��#�x�hn=D���\a4�N\Xx,����Z&�gyH����V��ڥз|��a$S�km�\���{^���q9�z*��s��
�V_��,��J��O���*p@- }�QM ��>�0Λ��~���5���K�y���+5{Hp�i�@qe�8�>t��5�K��M�}P${_swqmL���3�֧N����e���5�����φ���� �o3P}�򗣚"`nV1�?oe�0��X���H�$�3����P�ߏJy��uG�\Ě+z#��V�������L"U�]vt+}=�LP0��c��Ps�T�0�v���rg��u�]	�B��IhG-��Xg��1��eՑLHd��Z�8Y�i��p?�ļ�'����ku���H2c�+�ų�45���'�C}�z���zVx�M�̭���7/��S"�،O� r1��{=(��&�HP<9]}+OR����<�Q��Z<�er���,Tv�5auIeE����)�R�4.U�,�m��e;�U��[t,[ZU%.���Nx���]8}5��~m」�J���P���p�H��)�Pw[6���f�h�tSn$3���vZs3fivk�*5S{wj�Yu�ax#O����{j�a�j�8oͺ�/1�O3�s���� �����ep=�^���� ^ ��c�r�f��-�&=oc��������o�� ˅e #�@U�j������V��ŮP�XݗX�ceǺ��	ξ�Ѿ����l�cN��M��>6.ց����C'mO#��P�� 6�[2�`�1]VL�X$�1���Q���J9d_�YPkĬȠP���U^���^�/L`��[������@Ê��Y�	]f� vit�lB�>�����Y\������l���-F*�m�
#`�/��+5\[o�[K�r��JI��Sۋ^�4��N1�J�hv��@� ����Ɩ�΀�u,+>E��.C�!�%V���WFJ9��[���B��1��T��0ki���9�8�c��lŬ�Т����Y��".�h�c@�|W#��e�s�o���)�{M)/ӂ�9T��p��I��R��m�kډ���!�y�t��] �?8A�rӁ�-R:�� �x�g����8��]{ ̺GL��)�{��:&�4všD��@���0v�sVhM�T�Ğ皀#ɡ��B����N�W ��?+A�fu,z�ۜ�j!��u���r��"�${ C3���;�J52�ZE�ҁa�T�X���$�&���Y���.�ՇY()C2~{���n����Vq.1p����B bc�t�Q e��J9k&0�
7��KC�A����7pI��n�/|���.�DꖗY�e�x�㯶%���%vƽ���N-�"�a��[ԍ(���r a(��1Ec ��1��c��]�E�u��]��¥��+�db�a�?�[*h���(+]�Po����J�ԡ����c\�Z+HF�NQMc���l4 ��D�J���)�fz��ꕱ2擺bimI��؉N��ܜ�������@*ġ{��xf���O"�31�:�惧\pt�0��Yܶ�V��ﲨܓ5��1��٪�'	��X 7
PU�Z�%r�zn���ۜ���D@#�7�A_��[�,���R�OV�R����_�B��qd��䑹�E�"����� O��׭is�Y�� �K^��FTv���k0�*����R�Y��D]���x�,���n�x�n�{r/W��1N����g=P����kV���`V�-wo�W�6Jڴ��mV��	 {��7#̋�q�	�n�gu~���ߘm�'˷���)�Y�p��rg��!�X�
�iu��}F����(6��wE�n��AC����:��?��ɫ��Adwr0٤��;�%�/z����"YK�w��$~r��� ��5�z��k5^�"C(��[9?�h��卬�(Jۏ)�N�<�sh�q�����uE%EaqY����cu7fq�>�[�n���vY/��\�A�L��Wj���+`z�1�z9�٨�UA+�Jtu(��~�D��.�EK$�z�a\fi�@z���eɖߩX�֒Ok�ulQS�����ރݍ���٠7l�A�sl�^f��,"d�oU/�/�r
 ��J�F=zwI��?a|~��3
(�.cjP�-�~���:Yʾ��"m��3_�@m�1�Tҧ�S��(`�j5Zv{�w�����J��i��n[�
j��M|��$!5��WA�g�Kb�c|�,��Μ肊0;�ź:Ȁ���j���}��	��)0B�/ ��$X'�>�z�]�.Bv��E�q�����f�Pd��ac�ن�-����O�@(������;���)����YR���F�zD� M��1�|>S�^���5R{1C�¢a�\�QB)l��.�얘XЁ���pux�ʆsګ�n7�zqd&J�OM�9�ڔy�6�SfV×��&״]c��$���Q䯬�b�]�c�8�^�v�q�z���r�ϟ
�]g�w�$��=����\�F��C�8D���w+�}��~*�$?ʠ@.A�{�ţ��v���m�)�,r��vsh)%_��u��}?H!0d�@�_��(+\�R�R���R$Ǆ�zG����Tw��+U��;9�4��+kNߌ��lY ���:��f�al҂"�Y-��vf���{���Le^,"��y���Eu�p7vW:&�L,��l!1��Q��YhB��m�K�I��g���6��?�k/��Y��[ito��U�®��1��l~-��.27�Y�r�=I�L��wn�e��u��(��/�O(�������*�o�C�]ۼ+Ə�-�*���#vz�R,�#�s�K�)+i�cZ[���b���b>�rBV�:��S{��c�l�$IԤF�����/��L���kPQ�z��~!�^�z�I�Օ0���������3e��d�S��e��CM������{��s�h
�K���	)6,������+�/��倵c��D��B�w�|e}�#ֈk_~,���om۲�'��ܬ��?ؓ�/f%>T�n�������	�
�]�mk���0h��v�m�Ϲdۻ��2��cB�#���R�?�Hj�"�r��Y2�?|D���y.�K(�ҁO2��+UTg�����d9gɹ$��z�6O��x�F�Xfjp�8�u(/�ůA��>y��(yЩ?�9w�T�N55@U�7yD۝�����f��,X�����pU�<+�i�%SQ�W�W���zII1凎�^z�<%�ɣT��֚��}�V���v�w�ѿH/�uL���ǰ�h�OC�_�${y}UCV�_�I�����Q� ��_s�,�Gq&�	9��SU� ����PCYzL^�؋��;>eυp"�ٽe�O[s�(���L�O�ó1�¡���4n�h�UvAa�1��*��$+��T��+�-�[��ؿ��F�xfT52>V7F����!��k����M�r�V'�:<���v��;2m���]_k��̸g�c�4<z���=IH��W��%;��h�Kl|O�t�#&2��B���_�-�L�O����z�FS3��	縌+���*�>�sQ1E!+�IdJ������bA6c��VG�B�Z� �Ƴ�µ�趱S�����So�	v,Y�s�
t�>n�+��Uk[f���rCj� �Z�_�I����{L5�V���K+q¾6j6H:r=�s!��ʂ!V�|��BI�6�����ś�� x/�ɖ�)�R�iH%�r��J٦hk�$�i�%��z�K������~	`�.3�pulloq�(?��Q�T^����x�'!�@B@�|nU��M�9������p>=�s{�^Pw����J�ɩ�%��{-�[���%���M���������}��qdJ�|�s�~��MM\�����͌�ܵi��Ղ'���R�J��uo[���@�l�P��Hq�1p� ȏ���!Ҵ
�h\n�,yN��;`�� ְ�s�	0�)�f\5�'B$��+~(E0�RYz���Yr�ԅ�
K�:���WF'����p^��m+g%)��G�����(��$m���bu�Y�a��Qǎ� �T�H��Żt^|O;]xC۲�S|�+OӖx��
ub`�aV�zmJ��庖Ϊ���P}`ć��5�L|���İ��4$��2㑀d�[E_.���B�����K	kTܖ�Y��-�2g�_#J��y�*i� �^�%o	9�uƈGu)����<�˱I55o���=�G�M��H�iT���:��PQD�
��/!��2��/�Q�ެm�A�>���1W6�A[�"�����g�G	dIT��B�{��cZp�3<B0H���`�g����y�E�ҿwv��V�^�a��Am���w.Q���e�&� �̨�{wK���w��{SP�s5�RW�
&R�'��q�L�����k���Ւ�V%G���ӎ~R+���z��+E<�݁�a�d���|t([�T�j
���F+�l=w�'���s�i7ζ��ߙ�a�DO?�rD���g䊘�[���7���M��>s�z�[޳�౦�_m]	v�Ѝ�L�Ì�C��0|/�	��P��/UN<�z�.kjΛ���8N<� =�xr�	.(��ֲ[8�Zs�\|n�X��pt�n�{F:�LT?٢+��Q�&9��
��ZX�h�O����S�OE"��P��W#�<nqRn�X�$�.��̆M�K/���|��\��k������{�b�v���V6�����&���!r�@��w$�
{a� ���e"juI�u�.Y+c��NZ2�� �M���A�2�1�)w� �ܫ�N�IZ���)��fU�㟿Yx+1��&���Q
,��pK�+*�>֏� r��0n�ak"Xk�^��!�5�(���}���q39�9�My��n�_�o�@y�cjʋ}pj՚�=�΍ܕ�d6�sЬǂRq6���z5O!S�����FD�9��r��EӻOa�g4|�ubv�SX��C!����W�&<?}t�]u�-+d[�[��&��Cn�������і��=QU"8��l!L����	���y���JQ5����#�qbn�Z�0)Y��1~� 3���ޮ̈/�sv�mт*f�1&iDݳ���ȓ�_}�|��<*ڵfݲ�.Ly�d�1Kn���Q ��0�7[XhƳaIZ���i���Ӽ�hMDZ�<�5D��[N�M$�Us�J�~r��:7M�u�����t���c�i��vҺ=��i��D� �1�sZZ�,�i}~�iP�鿶F�N�e ���O�t��b+�kI�����f�LJ贡E`܉%E��#���=qFᑘ�|}��Ց��[�<gYZ�1��"B��|���LG�<M�Rq��@4�4I�_�%r��	��.�\&�	4�-^�����P�"�Q�ϕ���Ze����f����8��Sb|������.�G��	��c-�E��9
Y���٤�d�;¿!-S�����C��y�v�F�8�c+ޅR��_x������)E�Y�w�5K�����"�V��C��>�(�	m�R⓶5[1��Ǉ�*�� �.�W#�а�H*���{B��5<��b��w� �s���P���	`�P�OyQο�b���}F�-����d�h|�p�P���]�v�`��`�d�|�
KN"�(�^�F�
P+�r���e�\Ś��������
���!�:zt���s [G��-�¯)WݎK|hC��Z�}�=�Bt�J���}[]I��^(���P6$z�Q*6��	��i��B�\ρ{ڏ?��ڪ�3��|Dk*������\�ߕ�r� �b�xq��Fs,<��C�� �uJSg���_��	���0,��^��Pݽ�A�۞���j����NHL�Ĭ�^=8'���̊&5Ԃݖ8�!{���t1[�~MH��\D�� ձa��h �S�@H�9]ċۄ�EkP ��5�ua̅/���n�^,��6A�U����J)���(�)��h������7 �)]�c?�����~�oS!�P+��1T1�:��,d��]^��-�O�j��l�E���?)��&"���2��ތd[�l�9%�&�T"�&��5�_��'�5�ʼI��w/-Ά�u{����K����7��ߔ/hp x�������{�D/�Μ
�#�x3��O`�h�R��-�0oF�=�{��d\��p^`�4�P	�I�@B�*r� }��f��6�e���d��ɖ���l����l���� ������˸�ߋR/�����q�2�.0jk�f�܊������a�Ǌ�ܬ�Z�����YTA�r���~�6G�oN*��j�ݞ��|x��:����ߔ���|Q�y]۶�<~��꒿"�X�А�
��}b݀��չ����+a�)&���9C�+V��Z��ht-<\J4��й}ǬW=C�Ō��6!�Q���v+]��з�5]��n�q�����#_�)��4ۄ��L�\���l{Q����[�*ZD��:2�V ��v8�c�ߩ�Gי�8�<N�����:|�{�5����^<TV
Ð��$߳��6%`�	�O��{�#i94`�`�ɣt��cDi�N�y��h��4�c�t"�m{�!*e�>#��������;�/�f���VѼ)N��(�e&F�����i��)+��x�+�U���$�z��2դ�?��
��ځ�h�,P��6��T�V���9��=�G��EΆ��+�q�DK\�e'��8����j���W���!l��}�Ƌ��8���&�ޯx��q���i��U�?�k �!����$�R�e#�r��5���-�� k$$,�7O	�kI.���4�^p\���s'����>=8=�����&&I�2��|�RQ�t��֢-����lC��Q[u�芯_���Ӈ��eU��� ��ϻ@�#���@��M^���Z�v9��_��
�i����78gP��&Rb�ĥ!��m��*,o$bL�ۼ�*����?�w.%/-9�%�e��e���%,$ڨ0�4����,C5vaP6�pp�bjT���ï3�$�@ߘ��/�m.!�OQ�T���ۭ���%ڴO�I*Q3�m��I��}8���#�PD)��т���������fנ[�۞���!����C�=�O�*�6��-2����>a��u/����b^�}d��WΌ�,wN`�&��-4�Z���
_�*��/թ}C����TI��Z���{.�RSߠ�
C9����$���Y_y�����Ȅ�W�F�^���+]R
�v� ����cj��<��H�<��Y����!��uR�6@�=��5��}�������ә��{7Yf�0۠��_@��%���۝=�5���{�����Ȭfz�O�˦�cM�����].Y�KNҨw����fm>�|�5n���ۼ��6<$�e.AҾ�d�ǣe#Ool���t���vr��6m;3L�sC��ڛ��Z�Ġ8q��L!&�KA��[ ��Qav��\��	�9	�Ǧcvc�-�Z߸z���R�ڧ��c$�W�(�`��,�T�R�vē)�3n��Zn�V I�gX�]� �F����<���,�+�EÃ�')�S �?����5�WvfX�_�Q:T�d�8�:0tL[�+��[u��/�߾d3[���o,14��o{�cF|�F�*�T���q�`B����z��Z�Wc��%�!%VA�g�|���3���	 y��i�Ъ(n��&݊;ؙ��I�z�#�R�䵪�_�Z��r�����_F���M{6�)S��=c�)�ƻz M�J_r(���L>-Z_�<�;a��x��l�C�D:V������$��`IŏQ�>�t��s��Q^_��7'׎$�y�kDi�l������$�`e�6�+̠����tD'fS� U�f���*:R��k�8�5�-tR�c0d�0�,�7�9�\ŜF��܇�5�9^9>�1*��Q'W"�c�+�Nvq���W$���"1|H��Q�˙�B��F�����5Ii�w��A��q`���f�2MԮ�W�vf�l43��Za�n�D��\"����&�5��[)�Q�+0㙘3����KW"u��ٍ��}E�&X�+��*��]�	t�p`P)=u�d��R\ ǵ�/.� L!A^{tog�#5���}��H�O\�H��-�1Ͽ2�F�wN�S͍������R"��� .\�i9T�F)AIc@��D�3��ݭ�ɗ���8喧��$g���41E��D�*"����OnŜh�B�g ����Y�i)wU���cZ,U��C��wlo�5@�<�e���ݣ&(��e�q�厄.n^��83��2(�� E����hn�������&*�E+�V�8�r�hv�����uKu��q�n0����.?����W]8����yI�!���	L�c��xu�x�1 +��-F����Q���n˰���ܿx`>f�#LG��n��e�m�PH���M�g�kI�.�S��W|n'#�F+�������F�o��R�rt��ˌ}�U�B��S��+̒4���9M>���{P,I��'��cF�C��s������i��<7��!�*�� r�!�.�"͚u����emB��+2��Y��֜�C��E��4Gp�
Qn��gH�uu ���`79L��q=t�������a�:�Bl����������l���9���6)��he.Vc�x�;�xˣK�-՟B|�d�B�S:�ڊ�-tw)�������#B�]}�u*55g�8�c����9-�n���Q���ѵ�Q ���������:�t*���'R�ZP�E�.��p
~���r�X;U&C���v���|���.�kq1����a����`^l�g �2��)P+�U4V ��b����'�\�u�A����>�:]N�B~�Q�2t?�of55wn���ʃ�G�����V��|*�� |����ٍ��M��H��ʷ�ް��[#��
[8��u�&�5:u8�'P�U(�J_�Y�O>'u
���E�Ց����P��#�� ������e�z�*�!0��7�����N�f�6aRy�w������0zޕ��\Ĵ�q5��yC��9T�#��<}�Q~�����X
//�$ �p�G����~{�{X�}�}Ko�)��%3L���Mt22�x�z�b4�l�D�# I<��+�fN�������^�������Kj8!�!>wKv�=2���ZJ�N�¨R��
A��l���u�_8
U4�O?X�B��$�l�9�����;���~�3����k�=E	��[�:`{��Tn\IM4�J1���#I�,����E2�ڏ������u�=��l����=b�}ۆ�!NV0�|�_RS#j�~��#5ϕa��DpצSQ��S�ү�NNa��h��gfb�~�yet�z}��t�-L7 ��[s���0�s�v�*>�TGϪ�@���`�X�B]q�|�8��7�׎��O����Px%ˆ��X__���Q�*�%�՝FK��%�d5u�_�馊�g�"�`�}z�6 7�$�\�Qo���tT0+WVК��~����b�1F�b�m'�Ɉ;�t
��Ke�8����2Dj���*�8#�Wh�!q��P�y`X�ϣoc���.��1�L*Q0�&�%�6�`�϶9�Txt�D({9k�y&v�]b/���DY�щn�۔TN�N���g�:p���:?�$VoEt�%D�s�b@���g�k���8�T$@�6��������d����Xb���t*�͞�x!�83���G�C{�T�s�Hü�o�c;1=Q}m::J}U�x��T�����Ώ�K�w)Z+�>��ʙ���l��t�&�Ou��i�r�?��1Wl�$}�C�)����,?�l��kq���)?'jhIƔ~5�����&�r ���\T��*��[��5IVv��{ l����Oa^�'֡屡�f2�x��t^���L�T*Ss��\�f��*_$;sI���N3�Mk��Rk�|R2�)价4�$��2�U}Ps����3&@Q�=i$m�8�活�����(�B�%6c�'� t�>,�Ϡ8^�0�L�	}<���� ����[��.-B{l���4�ܖ�7$�v-Y"ɪK��wi��A(�u���©`��k�7+����8j�;���;b��I�qWUA��;f���Q���y�29�p�=�D����y�����է�o��\�غ��f�IT�U-���j�#V��or _���kTW4n[%�A�&Z���������m�"����Q�(���/��Y@V��a�'s^'�br�ǧ�O߀X`�t�B_mW-(O"%~lIr�S����y:����z���Mzx���,��@BQ\l���k�i\�� ��+�$�(hM2{W({�&��jAP�F���rp��i�w�\Zf��f��E?�I�a��+`5M�V�1i����7��^;T$��O޼�_'3��/R�}ڏE|<�o���`�i�'=���A�o�`E���e4�9r�s�ۍ~��x�0�����Q��������n��k9-�R2���/=��+U�C�h��`gZ��r��GC&( )6.d6�_���?t��J�Ib�o��%ς�>��*y}�s�=ʡ��~=X��X��_��ԱȅU4�d��Z�^�cѽ*e[w੩}��4�T�2A|G�%���M��[�uʷ�3\��Rb:���d&�Ye�����;���ϤO��.jm�yx�C�0FH��m�z�˒PDM��Ktl���gG��e�_��m6���\f��o%�uR7�n*A�9"ͮA� �w-�C��]��=�竊sK�?�6z���)�4�b�=�mP���<�D@	���Z��t5?U�^��'���n�d���ؠAk���~9�#�j6��Tj0_&U<�C���R������A늎pv7��O�N��)������u��x������
���r�=�#�\;t̗���J�������y���bG�>}�	#H�尳���v�&OU$c�u1��\+�鼿E��̌z�!K%�&��������Ll�/Ja�RB7uNTeG����p��	c�a�B�g�"b���w������ϲT�w/)6C���mp)�).W$��-�B|C�>��8�S��z���u->�R��r�W�"nh�ɔ ?G�+#|V��׿k�<�os��'h�&����wh���JZ�w��W��}>RbNwe�Q|�eYS|YY�����6�`��OJ���q���4J�4"�zzlކ�P�ƅw*���|1��qۗ \�c�5�eҹ;�� ��Ug��q������ۓ�sD;z�U'����礦BL25gZ�G�E�?��B�K��їZ}�9��Z��L��۲r�Zi川n����8HZ����SN9
�U��*����Q__���������~~S"l��r\Oa�i���XˎY�.����u16g4��6l�%[5�݂i�+O�6��,D�3��[�=oo(I������?���5n�.I�u��pi�o\���2�􄸇��t[G���IJ������X�M�E��SEbV�^��O�h/S;��trK� �~=�)�u7ҵL�č?� �D*w��Z�������
Ҹk�B�օ�3����巧xvwܕ6!��Ż�ΆX]m+��tqv�e�M9��ڳzP�O���f@P��;s�e��JA0ܞډ�||?Zc"7��nn��p�OXkm�r�
]Yi��qLcڲ�k�@�V��i��?3#�zG7����Bp����+�����Qm�E�'�n�9-ˁX{2�������^^'f%�����\���,���k��Ӣ��[��Ir#9Y�T6���"����HnH;7Y��SX��R�9C�`M	/����W�08[�Z�5��YK���d�il��Y�����/���E�<�6��a=I���=��'�]�moH�-��!��]�IX��%"V_m�:̢3��G��S���{G�.Q4�N5�|_\Ё5���ґI&s��b�����\Q���U�b�M��!:�j�ށ3�-��u�=�����3���+ղhm�X�99�8�)�;e�"��2g�����@��+:
�s�f{����ޥ 8ZU[��3J��bs9��3�ME6��<��<�UnBwi�zv�Z?�E`#��ޠ��?*s��SM��G��W�?�|+�e��<]����"܄��.܃Z���$�3��l#~ũ!'SK΁�mnOAL��)W�Ԛ�a��<�p�W���ߺR_H�Mˇ�@)���ޭ�����8���R\?k:`��S��"���T��Ch;n'����a!^��l�'��?�FǤ+8�ҧ�t^I�=���s�D�G6O����;�	��$ƻ�CNG�V�s�F��)�_�a�L�����?M;��V�	zC�~�g��]=މ��f=�J�X'P˽�&Kj�e���/yO���}F��ͅ
��vT�W[IϤ١w�'�sokm2����u��,��!6~�	>zmg���UVܑ�6�1�>ѱA�Ȭr(��'�'�@9���oQI"�d͞?�M�b�1�*z^��:��8��)�E�M�p�4��c�!�u�qݞS�-��&�xl[�5�'�^��?��qΏr�Aq�	�b� u�月��$�{�!�L�J|8�>kCMN��k�dH@E�
�lDɈ�y�x	DcCZBDV�����VS�+ioQ��������8���^L4�(My�L< Ǯ�V����&R�9�sOL��/mM�5.Ӊ����(�]�d�A��������]�d˶v�4�ʂ�@ٰ�C1#1܈�]r�/�U������*�3��T�w����QG3�M�(5�=��3$�E��[�P|!v�4����0X���q�&��|9���kf�W�Leꩽ� �{�~<R!���ci�zO�G��$Rn�7����Bc%
�AzZy�����>w��Ye�D�]�Ǜ�|U���g�������P��t����,�E-��K���'iIوC�$C����Ks���@L`�4j��h��.$c��z�V�,�կX����B�)��U�6YM�I�^+kQ ��a� ��ߠ���х��R�k)���,���We�
oi	y�m�?5�V�W�V��,�\ ��w�6����LGQ&�x7p\QH��z��8�}����R���G@&���O���`@=+��Į��3�'Q�C���ҾuWxqp\����M��˺��{nR5ʐ�Q;{-g��?-"��\��VT�|q�H��Ӗ��(tB*��^bZhEۙ�wL`c�Z�(���#�
M��Ys�`}Z5�I@i�tܪ�;ח��Z��!�ԿH$<>��Ǔ�m���� �����Sr)���sA�w��t������mUmvTsZf��}ԥ���E��Z�XL����S��Z�����E<,�da'�6-x����|���.E-��a߽��-}�s����1,0�A�2�"�	��tq�<����c��5�։�~���l�U$D���m�0��zɨV�t�� Lǣ���(jޫ�(m�$QZ2�8���_���X�0��ѝ��4W���v[}P.΄?��6��"a��U��U�~��E�Ӭ<i(Q�gNp�t�wi	�0#	��֣Dd�#[�;�@�a��W����m^<ZX�(�����3y�~�	�C��U�N$��.����� t��;d�jvH�pGg���d���Z�{9�~]>��$T� s�K�50ӭĸm\�P�ҍ��j������O� ���~_��]'y�X\���$��jqNx�ҷ�=OG�a�G5��j�a �y�C�/��)"���]٬+%����qB���2��V��r�y�D�	������h#��A�@��Qq^�ز�&�������}�ƃ��K����غ�ճ��T�"���X_��ܫQƋm�7� ���"��/�p��1�8v�X{����<B��a^�T`�P^��؊A���%�r\��ٺ�=������Go���6єsH���Q�ig&���p��r�X	�<����.��Y;�p�^k�B��������m�'ё�� �ᘷ}v��\tx+�ؑ��i�{	Q� ������dpFm�o�������%�-[�o��MUw�O¶�ϚAC�H����膈��e�y���phn������u�W7󯅻$��56�8��	̩��X/Т�5W4C��`�'����o�<2D���x���#��lҔ"��s4�g�Ms�np�s�?�j,F ٪�ҁ^�a�1l߄B=
y�k��'p:VǙ;>�H<�H3&2�����z��sN�E��Dc�����c~�χz������GYOL\�	[t�*���ӟ�~��O� ��A]+ɿ�$�Y��XAc����Z�.�I�%�L��Z�Ԧ��������<l�Gu�$��ԙNV���T��t=�����ڽg��\���!2���b���ww���2��L�|�h}��� M)m��l�,cN!�0iYIӹq�H�aʚ�����w�Q�3��<�T�R�V��M�������U�J�\�����+�-����N�N�U�b	2Ɋ�����	���t():.�:����0��ݢ"��M��im���ص$�{(x���#��CE�<���2w��d�|��[g��Y�R�^��	_������K� ��3����L�l1W�m0˹�<�eY3ڟ�3c/��Q|#[�;(��� �˽��`$@)��9P�A�P�C��)yj�u��*+��D� �̒2$tgi�Myۢ�����{���%��(��Y&}�ZN�\0�����;��v�?��1���E������ƫ<-�o�9[�0n9�<{WӞ�Ӻ[��蕆Ȕ=M������M������R2�=����S4���Uk�Am��i$�9bWBU�mm���t�O/�mcL'���V�	����h`Kr��d
�fП���(s�
Χ��j&��zp��k%���nt�Ϯ���j��z��?�J��F	0���>�
~�Wh"G�Յ��<��K�~����
Ƌ=��w���~�oϑc��8��&�����ϡ�Ծ��K7?�@�9��#�� ����y��ApNk,�2��*=�����<���dԻv���{�qDX��z�%{�(g�D<7l��鸆���h+�c����.\���P�)~܎��X�3���^��v�+r���,%�T��6���^�%��%�%kE�C�[����k_ˋ��iV����	���>�/]�M�D�pA����X��Ӑ�@��8��A�����4�Y�7t�E��E�ǯ񓧢I�����bI�-櫚�UZ�b��n�d;�x�6�=�TA[�Z�E���;��>�+�}Q�u�sG>�?v���
ѧi(7�}7.������)+�4��P��Ȯ>+�a������c$I��D�4��aL�6s�D����4#r»�I�����-,Y���ɡ)Ϣ�>ڇ�5/Y�{��U��t���q1z�yH�����6~�R�k��0�����H�@�N�ٗQ6ܑ���v����ļ�Q�4�eTD�>�tYN�S�&��v@��,��\P���|x�{�0����7\�z��{�r��U�É�Ќ��\T�"%�ͩ�4�OCо�^)&�~�
F�])m�����hڋ%B9�vzd8JQ.V0m�������j�Ă.���ɏe�՜c]c�7��4�aDWO��k�9�*�:�Q}�O�o˵��|~�pai�N�%6�J�~�
n=�9�R���f�V˄\}���f��6W�	=F͂�0�` ?�|\���t������,�sF�V�F��z^��H��@oXKb�cE�!VM�%d,)���1�B?1y:! �ڪ<�Pi���G��u�������Zn*
/Uf�H;E�G�B|1�3tU(��X_]
��gJޓ�Ts�,4��Iȹ���g<���pSJ��hD��x�v�H�ëA��Nˍp[Aw�gq�����7k	�6�c�*>\��i|�o�:*�(X��c�$����?��oP��e�˦\4�|�!��`V��h@���}�4��슗z�K����bf����Sb[�V�Ũ Y��L��v4M��SV͸��7����(��AJ���b�0?�'��+ cd��Gҁ����;��@=R���4<-a���hj�֥�?�:�-�ۇB��1�2�,���	����j�z,+��e�P,1�&{�&eSUZP�nĆ��!�Z��9暾�4.\;1.�r Ԋ0e!��{��;�8���R_TG�������#��I����Sٴ�3g�0��Ų֢fꊨ'ڽx�a���R��(��٫�6.�T8fE�rr(Ï�>�&�Z#"���&0����KS�M��h>2/ζ�&�"s�t�0�>r,V��`�l�� ��T���邋 ����.�j��`�`�o?�mCj[�i'��<X�ޤ�<,��8'P�(����}��!�o��ͤ�e�D����y> �`��[	�����ǡ��8� �L��9�ʢD���r8O{�	R&�B��L��{Ɛ�j�B��w�c��#��ö�&ۢ��U6�T�6�w.샇w[nB���r=azywٕ�K>��Q�UMG��t�ܩwXa(N.��{ý�e���w��9�?�����1�svv<r�
ؚ�]_<�=�PT0���g��v �JG<i�]�a��MB�X�	�Av]��''�0B������/f��q����������zmSt+B^n%u���q�j�lt;H���oy[���1zS�^���M��.q���LVĥ�L�9 ~��Ѯ��u������PA�I��Q0	דV@f\`}��9��������;�~�	t�1�S>&!.4X1c;�6����Y^}��Pz��z(�����-��C�0�`��qӥ�B^\�'�cleb��Į���}eIݣM���U̒އ�Є%6��	����d��u-4�Tp�Oq�џ"0OR��5�9s�#�<���j�V��g���"�GIp�n�e�י���k�@�0c�bl�k �U��Q|�+����CVğ�]ǜ$%�} �&��Kxm�<@�<�|s�}
����0
`wP!sp��Wx������X�'��'�¿U�#��>pi�R�b�G+���6<���������fO4�u�]�l���}��bӟ��r6T��w��a�5p�.�O�.F��uɰ�g���1'��6��4����(b�����|x�#Yh�ְa�2�q�O��j�-����Ǳj��?�j���\��4~G�$2�.�t@�#O���=d�o,���;Eaﰭ��+���.(��y�,�����cC9$>���ϯ��c�i�m���@�p�%�!<l�G��ν���Ař�J�w:�!{i��@L@�'�������e-�J�Z�')x�?7��u���^B�t������sV��6˝ci�-�|�й{�3>8����ʳ,-��!�����0��:�6�T��S��og	���YQ��k��Z��V��_D>��^M������v�s�~cL�*�AI�oz�جB��"�׹���?��zf�EO�?F�a@�ޟN�YST�����,�ʟ��f�B~�l�XEj��Yv�%_;�S��zV�(�1>�D�/�!�!윜U�Ϩ7�ݗ�,wx��e����3qs�c<s�	�Ǆq�Yح	�ذ�F]1]T#�X���b�P6�'Ѿ�Z�{-��2�E�ށb3�>����6��!UOK�i�e���*�L(���w -6�G�:;Ί<���M�`8oi���sn�Y���b��{�"��:��AS�v��>qh7�7�Lni�5 ����V�	��bt���fZ����r2G2s���Hy����e�<�,��=��q�]�R�U���z�Қ�&�7��k��C��i�n[&��h
��2l^�jNj͵�>���\=) @� [i�OɆHҦ|:e�x�[arh��x��;c�]PK`�K �U�< ����%�XK2Ƙf��i����q�-����@-u�@ 
�	�L(G �ة)�;��a���:�{�V�[N0!z�z�伞�~R/b��;�[��8�i�Ol@1}^��*�<�-8�PZf��z��>Q�ܰ	EI{񻁲'-�kt�+��,�g�h#BV����5��U���d��n ��̙�g��l�-FԂ������F��XG)d� �R�Fȴ��{L�,"��Q�(
Ұw��}��q�K�,�1�����]Np\u�$�z���d�0ɵ�)�Ά%|�Nb.�
H\��:�;����G-�1�>/�'����T�c��xi0�RSb :��0Z-���\�΀�|z4�t�9��61���}}�Ƨ�q�$ӿ�5��2^W����cp5�R�x�^\�>�����mx�1I��:�j��� �s��x��%����=b���j7��\isҡ	AT�~����Cu�g���k�4�P�7���'9#���ӞR�B��1���ΛkL\[�k��4ӑ::���}k�U���^Ѓ�]r�!�5b�w\��!�b7��Y��v�����©=�¦�ӱ�,9��=�g���~�����8����d�+ĩ)�b{^��H���Y��T�$�2F�m6�ed��9�g=�o�>���2���\�խ���{-�X��B��uԵz\���Z�rˊK�MA�r��qZ �h���@��r	�,0֒���&(�zmd&�����t8-쇁;wɍXc|�N�� C��Qn�vP6����m)�`90��^�N�b�br�F��R�5ݳ�u!�`��HѨ)��:2�)\t����㣓�ɞX�'�3��࠵eL��/�$h'3�R?�f�`X����kg�2���U�F��ߊ%�^f����mCV5��$h�����n��$[@+� �e5�lfI���.JR�s�sJ<���热��	���c-%�����o����@�����8h�w2��o�9��;lO?�d�T��#
xx�}U��^��k*��3��eUB�1���/~D-B��S��Pc���(�J���Ft��>_�n,��Lg�8o@�I�h�.���R���M �B�}�����O-��
z�yLw.�%��Vcj�Q[iAGe���Dǳ�-��:f�����l����:A�%߱~�OR
<M�7��-��P"Iy#�\�G����b��r*�}aSut�$$X��>Nv��)vv���c� @��qZ�B�<�@y�Jm�T����U���3 �Y?� ����%m���M��]�H�N~&�����w��\+e��3�4jHц�}��rxTTt����Ǩ�t�P�~� .���3 y
ΏA>Ǉ۞_�۾S���@?t�y=l�T�
����6�+>���J�_
�#���m��Jr����4�<ދ�T��K�Kc�^�[V�7�.��_+~�jݳ	��4�5�����n��a�pp�=�c
��@����Ϙ�1����_��\�(��[�Ӹ)��~�G�ެ�TS�ɑ|}�#L� \��x��sI�DZ58)��i�����R}j�4+i�Ok�Ki*�r�}a~�r�?���z��Js�]��%~@7Թ{��}P�1n��B�_ ����	M�W!<v����{Lʸ���e�9�c|k��Xв�dC�q�h��p*X�&B>�"G<�J�N�����.aIڵ�I���1$Ǻ���JF6&ŁD��$D��qwsbT��}����]l]T����f��f��G�)���4�` P?k\w����a.#����7�����t�8@�׹�g�F��,?�{�6�C�;�tݵ���r88w�ϊ����2)����
)�" Y �P�}o�%�0g�o
���'42�j�'%*�Wl�����
*%2��e>%�����]uCa�:�)�h�e�Z6��U�T(��Y�=��E���p��$�A<_�I�(��2���MX��
/��mS+M�Z�ˁ	����
m��6AӺ�՗s#�H�����'�^e�D���+󶙱��
|��Pw"»Y�)G�	*���<k�~pH�\X×b���ն��q9j�W	Q�lRB\?���t���,Ő;3&T�h�����X#�hXN��lr�^%O���@m��F2ȃ)V���i�<5���%柙�"l��v/�G�ү��Z�$�_/=�iN�9
qqy���^�u\������i	��e.n��,�y��d�~�Q�?����EGZ���݌�&���V5x���e�}(�_�}�[O:���,�[V\2�W�f�R�+,5�V;�x��F�D�`01����Q�J;c&�D�������X��9o�t�a��4��SY����e�%���7��*K��
�Q�&}��C=wF~�l�੥+�B`�N9�f����O��8J�y��E��iVf�e��	;�&mٖ�X�"0'���9Rc�p�C)�ƒZ�g*��'�� ��s��\`?`fd3_ZI纏�W�L��iT�#&aqw�Ox�<8����s\�w�?8�Ӂ]�D��c�Ct��{c?|��<�� ���Y������U�H�+d�AMf/zͩe�6G������[��͍���؈���p��B�.
ic�@ԇ0�����iyAF:7̏��A�(��He4/������T'MɜU��>���P/G��������-#7oj4)���אD�y�����hoT�w���% ���a�ݢiI"��W1�� c;m�8��h?��� t
�� ��lƼ�9���W5��U;��.n����	��w��q���;�������f!���	k��O�i
c
�q���?��T��2�K��(�q����}z�>��ޕU��I�u����	��Eh9t����@�IGjĄ�-�`8�;;PU�� ə3��1�t浽�]�y&��)O�.� ����붱� ¦3�d���֌��I����@�V��r��qh�������������=��i��!�p:���~��Ӳ���]G��俿zP-��,��\�2~��Gk���
^{n�u6@?#�σ�U�s�@���@.]ر˄��������3�
`�4�qa�ô	߲jm|�#�a��\����o@{��w<{J&w�JC7�Z���-�)	F���&����s���Kl���i3��lF�:Z0}�:��4
�m	��(G��H.CYe��Y?�8�p�y긼|�5^���X0Le��[�z����v�#N���� W�)Lm$���s�Mh芩�0�4eJ��)���"�D�]԰��&�8M�dhfi݈3:�1x�p�2˳⁞�	m{oӛ˓�K������ޘ�f\�zD�����CtaO'�U�/�7��8�	����1 �ed7a��(�[!��@Jt-�)}ջ\�&��Z�9N+eD���%�� ���6$����&6lW��������81���T��2�d��� Lt����׳�6]D�Obgq����Z��:<W���7-�i�H�cbi���3��=;;�b����<+O�;�(�>Cs䓀��ݧ{�l
5k��If�s�d+���ɣs9�C���K����q�|0�T����g����,�F e|,�64���i4��\�����#)R��D�����$е��J6z-�(ay��;��p�g<+g�h��S��$�wz�H���b�;� Krzߔ���>�- ������> \�p{:�*g�mgl}Uca!��V��I  k����}򝔜K�T$��O�����`�~�:EX��|������FH*��iA���n܀W.��4J�ys�\�w�c�+;^�QVX-a�ڜ��S���d��'[��ֶv�v^�F�U0����M��=!_�����$�Ԙ��跍�;:�:꺬�����$4H�F�D+��L=��>A����d��F���0?�-�N.V��Y,�45�����K��M������E$�t��	꺭k@D%���z�����M$:��]ط�X��<.$��\J1�0�a[��M�JS.�l�S�'��� ���P��+��O���}��@��x)����KL�I��y��9�e��"�m��;H�FT�͂�~���JsЧ�'�܃J&QȬv�C��v;S$/��s?n�ov�QC��(�1��q���Y�2i8d�(d���C\�"6�\�?� r����=��ۂF��?h�7cB��01�$|��G�#�ӚfyƄs���}�s&;2��k�.k��Z�Ik&�Z k��Ǻ�����$^6k7'�t��W̹Ja�(iR�^Aq�ɹڂQF�8n��u�	�@���igo��;��+U5�o� ��\h��`{��o:���]�:.N��ZÊ�Gz)�x�80�!s�mR	e9g��O�� �����`ۏ[�ǹB.����+v!��d�� ����f�����xދ0��4�~�˺ �������͢ ���G�b������T�\�
��%�zh�p���n��)h]���:O�\!&����5��06�ae�"��RGi�3j!�6��;>�j�8��D�Ҭ&}�ڼ��/#_H�u�O�[�"�Ȉ;=e1ކ5X�ƜI��_���^ ���W��x�]�,��Y�;��K�M�
>��<F�����[�B$�,,|��$;1s�g��Ui��ksQ�/�NY�=9�+�w�p������s�{�Q�#.�g�������F;���q��7�e �o E�{9��s���m���9t��y��[?H��nA����OP�_Su�:9pc&��`e��U����=W�6���Ny�o�W�vB@�\a���� ]_�9+'"p�ؙ.H��%�p�A�\,1b���)3�M+��aZS��`��x�I��d";~_?��*a�ne��	��EV�!���p�=1굏'�v�"���z�l�@��0��(ﮃ�{Oy��k�����G���3.�m�"�;(�	0c�8�HW�~��g���;>��5U������cH^�#:*��<�ԀE�Tz.��%:����=�`�Z����fo3�e�g�}��cKn��Ϣ����t���H��r?	�ԉ�0�p&x��GK���A;�	}bp�X�I'�~8�Li3ѣ�	8�r�M�iK�,Ɠ��y�j�20wܣ�����5��t0H�፮yR�Z��3�⩳M���Ԍ�O H2�L�k���WX#��2��M� H�I��e���^f6ו�~- ������Y���%X1��Z��B՞�����#�u��AT}j�m��]�kK��_ո�<2_u��PbSH�Y8�4�����������{?T��Vslrփ��i��G�&�U?�� �GY���%�#�M��9SM��Ðs��h
���U��W��i��МQ�̬v�E��q9�M"P����D;uya����~�I+	����/DR�߾�D����uzc*����F\tf�N+ꇘ\�2һ_�[����P��iT��j�����><�k��ڕ��oo��%(�p�a��
���_LA�Y���V7��B��,�*h��y&��;LE�G�y���7.pc�Z�r�F2?�o@Wa$��C�=��ݜ8��B*v����<$�����;�^C��{�|���t�Xl���4�Yn�TՆ��No���>�ٌ&�k~�R)��x�F��ݾf�o��r���oV����AUO��������	~��6�l����5D�n�Fh��0p�)[Sc �s���8�q������:��Ϊ�?�b�����b�©4���Ƒ�W�<�?|�������'8����B��XGG� (������[o���S���'������I��f�qV��|��,��,<�"��D$�|��t�É.kQ��4TP`�\�"�ScNE��5�N�Lt��ø�b"�75g#�S{��z���l|(���B���"��~4�8A��k_$�Fo|��y E �φ!��e��='����X]^?�DR��u���J�r�:���%�I:yi�������k��߿2���B���s��MqzCY�n��O|�t���8���݈��G� ���KF
٦��83�o����5�p�xz�Z���2 ��Y��L�s#����a��X�?)��x��
���S�޺�ed��ms�f�\5�e�qvKrI��}�72�	���j/4۾�ybUo-1y)����������&�ۧQ��qa�A���)f{Mg��:� E�TY^��f�y�	k����4�)�a���5�������ԢGvQ̚�	t+ ��j��,�̎�H�����%he̅�_^�g��6a�"$�T� ��!��k���$a+� � 4	�kB�H��j��EXWC�\E���*��{�-��� As�G<�A]ɷ04q��h�,���;�&���9�v���*���
s?��:B���i��
�s&��[���Zge<zYޫ%� _�7�I�t�}IH�ph;^c'͗�3�V�k�$o�p]I[E^xj�97(b�|I"�����$���5��p��C��A/�ĸ{�b:�V%���N!�GX�я�"���Wem+;)T����W�F8�i(B�CP�����?�
�I��ц�@0�ae��j' �u�lB�*��e u���L^.�S�2������ ���w���U�K����W1�~��E�O�\�h�I�����[�%c:B�<�K�P��L$���8�Wn��=�����zl�;��@=�u�֗���V�����I���ѲZ����ֺ1{���PǕ�k��F�65���h��NV�⤍�/�����-a�7�j+�Qn93W%��
4��ԏ�oR���/�h`qD��͐��>d�-��s3ox��D���L����z�X�ƃ�@��ea�+��$�h�YK��Ή��^��3� �:;���v�R�?C��*����Z�!A�����j,���K9�&s�ͺ�j!d����0�Е��JP͡7��A�_(����]�zɜ� �t�1^7.�<�&g��
覛Ru�܁��F�a�3��K��gX����1����oKݽg'1�0�^4�D�BJ	�i����DM�c��������]�.#c����e����٭L��n���h�ȡ���=+VP?�ަLK�Vw,��h�K�Eu����
ͥ���W�)��҃��9�������H~��r�7�==��唪�m�xyP��7>Ґ(�W�ѳ���e�>�I��2����x.I�\=�651鵦�5�$���\�����E���ȴ ��1]�t��O>���g��r��_����TK
����H�NE��A��^t��^9�pWT6�"���g�,��b:}�Bx����{��(�J�E���f a�A�"�\�/�;T�_g�<��./FG���N؊,�R@�Ԩ��:�q�M.0gJ�/�ʹ�;$�r��tȆMw�>� e
�+��|�L��:rwF���jqXrYpc���<��W!xN����?�;���C�������qr-��B<�x����L[p���=��6W�����km'���Bco��v�)J��@�Ył�1�_���q6��Rt�n^�O�ç"I�WC�۹U�QZ�y��łD����b13X����p���0�k�f�g9�
��,�iw���-BU �\�@�ϥ���h�ën�
]�јYj.�+�q.f(�����K�簬9+�źǃ��,-�.�D�!Fܼ�ܸp��� 7O�I�
�`Ȇ��Y��G�M�e�=蹚_�aݳ�+���ɰKu׽A^�grPF^�]���F�}�r"�@��?����H,,S|���'�*;��
a�v�2��OYs���zZmt@���_U"���'�d�#�/���`	�@㑗'�T<
39��ǨmSp���,���97*����q��悴[�_�8&��{�뫦&-��z��gn���� v�ym����"�ků�h-�Itc�q
4`nPRXb]69�$����5�ACAp�X�z
�κG2BJTo������Eĉ�(B��'���J�!�"�
W��#L���mRP�����j�?x��#���	cu�(�Ԗ)�2��	�{��F��
%�VKk�.aU�E�?������*I�{���ߎ)�粧��O�-I˼oMV�j ��)N'pR���+/]I�!�D1��U�Q�r���D��@>!0���9:t�@7QH2� ���0���\��M�T{��O�v��h�!�}�T��&E/By��5a�k�����ڑ�~�pyFM�g4�UX�"����h@>�u�mNSo�!*�&%E]/�*�(�$��"G�Z�Y`���Yo$��R��*���R������A�����ՠ��u3�(�E-�)� �w\�>�������#�B�d=a��g�퓢����ڝ���O��� ���t�U�nNYNM���P[��!�ǼJ/eٳ)rtZ�mA�#��L��胢_tT�wB<��~�dt�3%�i�c3L�u0�RN �-�6.#���3���L$���.�	�Ə������A�;O$��Ǻd�;�O�E�4_ �Nٺ�4d�e|�����[�	�z�zm0��}R���ל����1���d�~��|�p	���ۍ[g�b<P��Ϡ�l)����=R���t���cI