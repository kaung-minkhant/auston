// DECA_Qsys.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module DECA_Qsys (
		input  wire        clk_clk,                                       //                                 clk.clk
		input  wire [2:0]  ddr3_status_external_connection_export,        //     ddr3_status_external_connection.export
		input  wire [1:0]  dipsw_pio_export,                              //                           dipsw_pio.export
		output wire [7:0]  led_pio_export,                                //                             led_pio.export
		input  wire        mem_if_ddr3_emif_pll_ref_clk_clk,              //        mem_if_ddr3_emif_pll_ref_clk.clk
		output wire        mem_if_ddr3_emif_pll_sharing_pll_mem_clk,      //        mem_if_ddr3_emif_pll_sharing.pll_mem_clk
		output wire        mem_if_ddr3_emif_pll_sharing_pll_write_clk,    //                                    .pll_write_clk
		output wire        mem_if_ddr3_emif_pll_sharing_pll_locked,       //                                    .pll_locked
		output wire        mem_if_ddr3_emif_pll_sharing_pll_capture0_clk, //                                    .pll_capture0_clk
		output wire        mem_if_ddr3_emif_pll_sharing_pll_capture1_clk, //                                    .pll_capture1_clk
		output wire        mem_if_ddr3_emif_status_local_init_done,       //             mem_if_ddr3_emif_status.local_init_done
		output wire        mem_if_ddr3_emif_status_local_cal_success,     //                                    .local_cal_success
		output wire        mem_if_ddr3_emif_status_local_cal_fail,        //                                    .local_cal_fail
		output wire [14:0] memory_mem_a,                                  //                              memory.mem_a
		output wire [2:0]  memory_mem_ba,                                 //                                    .mem_ba
		inout  wire [0:0]  memory_mem_ck,                                 //                                    .mem_ck
		inout  wire [0:0]  memory_mem_ck_n,                               //                                    .mem_ck_n
		output wire [0:0]  memory_mem_cke,                                //                                    .mem_cke
		output wire [0:0]  memory_mem_cs_n,                               //                                    .mem_cs_n
		output wire [1:0]  memory_mem_dm,                                 //                                    .mem_dm
		output wire [0:0]  memory_mem_ras_n,                              //                                    .mem_ras_n
		output wire [0:0]  memory_mem_cas_n,                              //                                    .mem_cas_n
		output wire [0:0]  memory_mem_we_n,                               //                                    .mem_we_n
		output wire        memory_mem_reset_n,                            //                                    .mem_reset_n
		inout  wire [15:0] memory_mem_dq,                                 //                                    .mem_dq
		inout  wire [1:0]  memory_mem_dqs,                                //                                    .mem_dqs
		inout  wire [1:0]  memory_mem_dqs_n,                              //                                    .mem_dqs_n
		output wire [0:0]  memory_mem_odt,                                //                                    .mem_odt
		output wire        nenet_reg_reset_export,                        //                     nenet_reg_reset.export
		input  wire        pll_areset_conduit_export,                     //                  pll_areset_conduit.export
		output wire        pll_locked_conduit_export,                     //                  pll_locked_conduit.export
		output wire        pll_phasedone_conduit_export,                  //               pll_phasedone_conduit.export
		input  wire        reset_reset_n,                                 //                               reset.reset_n
		output wire        tse_mac_mac_mdio_connection_mdc,               //         tse_mac_mac_mdio_connection.mdc
		input  wire        tse_mac_mac_mdio_connection_mdio_in,           //                                    .mdio_in
		output wire        tse_mac_mac_mdio_connection_mdio_out,          //                                    .mdio_out
		output wire        tse_mac_mac_mdio_connection_mdio_oen,          //                                    .mdio_oen
		input  wire [3:0]  tse_mac_mac_mii_connection_mii_rx_d,           //          tse_mac_mac_mii_connection.mii_rx_d
		input  wire        tse_mac_mac_mii_connection_mii_rx_dv,          //                                    .mii_rx_dv
		input  wire        tse_mac_mac_mii_connection_mii_rx_err,         //                                    .mii_rx_err
		output wire [3:0]  tse_mac_mac_mii_connection_mii_tx_d,           //                                    .mii_tx_d
		output wire        tse_mac_mac_mii_connection_mii_tx_en,          //                                    .mii_tx_en
		output wire        tse_mac_mac_mii_connection_mii_tx_err,         //                                    .mii_tx_err
		input  wire        tse_mac_mac_mii_connection_mii_crs,            //                                    .mii_crs
		input  wire        tse_mac_mac_mii_connection_mii_col,            //                                    .mii_col
		input  wire        tse_mac_mac_misc_connection_ff_tx_crc_fwd,     //         tse_mac_mac_misc_connection.ff_tx_crc_fwd
		output wire        tse_mac_mac_misc_connection_ff_tx_septy,       //                                    .ff_tx_septy
		output wire        tse_mac_mac_misc_connection_tx_ff_uflow,       //                                    .tx_ff_uflow
		output wire        tse_mac_mac_misc_connection_ff_tx_a_full,      //                                    .ff_tx_a_full
		output wire        tse_mac_mac_misc_connection_ff_tx_a_empty,     //                                    .ff_tx_a_empty
		output wire [17:0] tse_mac_mac_misc_connection_rx_err_stat,       //                                    .rx_err_stat
		output wire [3:0]  tse_mac_mac_misc_connection_rx_frm_type,       //                                    .rx_frm_type
		output wire        tse_mac_mac_misc_connection_ff_rx_dsav,        //                                    .ff_rx_dsav
		output wire        tse_mac_mac_misc_connection_ff_rx_a_full,      //                                    .ff_rx_a_full
		output wire        tse_mac_mac_misc_connection_ff_rx_a_empty,     //                                    .ff_rx_a_empty
		input  wire        tse_mac_mac_status_connection_set_10,          //       tse_mac_mac_status_connection.set_10
		input  wire        tse_mac_mac_status_connection_set_1000,        //                                    .set_1000
		output wire        tse_mac_mac_status_connection_eth_mode,        //                                    .eth_mode
		output wire        tse_mac_mac_status_connection_ena_10,          //                                    .ena_10
		input  wire        tse_mac_pcs_mac_rx_clock_connection_clk,       // tse_mac_pcs_mac_rx_clock_connection.clk
		input  wire        tse_mac_pcs_mac_tx_clock_connection_clk,       // tse_mac_pcs_mac_tx_clock_connection.clk
		input  wire        user_pio_pushbtn_export                        //                    user_pio_pushbtn.export
	);

	wire         sgdma_tx_out_valid;                                                // sgdma_tx:out_valid -> tse_mac:ff_tx_wren
	wire  [31:0] sgdma_tx_out_data;                                                 // sgdma_tx:out_data -> tse_mac:ff_tx_data
	wire         sgdma_tx_out_ready;                                                // tse_mac:ff_tx_rdy -> sgdma_tx:out_ready
	wire         sgdma_tx_out_startofpacket;                                        // sgdma_tx:out_startofpacket -> tse_mac:ff_tx_sop
	wire         sgdma_tx_out_endofpacket;                                          // sgdma_tx:out_endofpacket -> tse_mac:ff_tx_eop
	wire         sgdma_tx_out_error;                                                // sgdma_tx:out_error -> tse_mac:ff_tx_err
	wire   [1:0] sgdma_tx_out_empty;                                                // sgdma_tx:out_empty -> tse_mac:ff_tx_mod
	wire         mem_if_ddr3_emif_afi_clk_clk;                                      // mem_if_ddr3_emif:afi_clk -> [mm_clock_crossing_bridge_0:m0_clk, mm_interconnect_2:mem_if_ddr3_emif_afi_clk_clk, rst_controller_005:clk]
	wire         pll_c0_clk;                                                        // pll:c0 -> [avalon_st_adapter:in_clk_0_clk, descriptor_memory:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, jtag_uart:clk, mm_clock_crossing_bridge_0:s0_clk, mm_interconnect_0:pll_c0_clk, mm_interconnect_1:pll_c0_clk, nios2_gen2:clk, rst_controller_001:clk, rst_controller_002:clk, sgdma_rx:clk, sgdma_tx:clk, slow_periph_bridge:s0_clk, tse_mac:clk, tse_mac:ff_rx_clk, tse_mac:ff_tx_clk]
	wire         pll_c2_clk;                                                        // pll:c2 -> [ddr3_status:clk, dipsw_pio:clk, high_res_timer:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, led_pio:clk, mm_interconnect_1:pll_c2_clk, nENET_reg_reset:clk, performance_counter:clk, rst_controller:clk, slow_periph_bridge:m0_clk, sys_timer:clk, sysid:clock, user_pio_pushbtn:clk]
	wire  [31:0] nios2_gen2_data_master_readdata;                                   // mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	wire         nios2_gen2_data_master_waitrequest;                                // mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	wire         nios2_gen2_data_master_debugaccess;                                // nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
	wire  [29:0] nios2_gen2_data_master_address;                                    // nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
	wire   [3:0] nios2_gen2_data_master_byteenable;                                 // nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
	wire         nios2_gen2_data_master_read;                                       // nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
	wire         nios2_gen2_data_master_readdatavalid;                              // mm_interconnect_0:nios2_gen2_data_master_readdatavalid -> nios2_gen2:d_readdatavalid
	wire         nios2_gen2_data_master_write;                                      // nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
	wire  [31:0] nios2_gen2_data_master_writedata;                                  // nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
	wire  [31:0] sgdma_rx_descriptor_read_readdata;                                 // mm_interconnect_0:sgdma_rx_descriptor_read_readdata -> sgdma_rx:descriptor_read_readdata
	wire         sgdma_rx_descriptor_read_waitrequest;                              // mm_interconnect_0:sgdma_rx_descriptor_read_waitrequest -> sgdma_rx:descriptor_read_waitrequest
	wire  [31:0] sgdma_rx_descriptor_read_address;                                  // sgdma_rx:descriptor_read_address -> mm_interconnect_0:sgdma_rx_descriptor_read_address
	wire         sgdma_rx_descriptor_read_read;                                     // sgdma_rx:descriptor_read_read -> mm_interconnect_0:sgdma_rx_descriptor_read_read
	wire         sgdma_rx_descriptor_read_readdatavalid;                            // mm_interconnect_0:sgdma_rx_descriptor_read_readdatavalid -> sgdma_rx:descriptor_read_readdatavalid
	wire  [31:0] sgdma_tx_descriptor_read_readdata;                                 // mm_interconnect_0:sgdma_tx_descriptor_read_readdata -> sgdma_tx:descriptor_read_readdata
	wire         sgdma_tx_descriptor_read_waitrequest;                              // mm_interconnect_0:sgdma_tx_descriptor_read_waitrequest -> sgdma_tx:descriptor_read_waitrequest
	wire  [31:0] sgdma_tx_descriptor_read_address;                                  // sgdma_tx:descriptor_read_address -> mm_interconnect_0:sgdma_tx_descriptor_read_address
	wire         sgdma_tx_descriptor_read_read;                                     // sgdma_tx:descriptor_read_read -> mm_interconnect_0:sgdma_tx_descriptor_read_read
	wire         sgdma_tx_descriptor_read_readdatavalid;                            // mm_interconnect_0:sgdma_tx_descriptor_read_readdatavalid -> sgdma_tx:descriptor_read_readdatavalid
	wire         sgdma_rx_descriptor_write_waitrequest;                             // mm_interconnect_0:sgdma_rx_descriptor_write_waitrequest -> sgdma_rx:descriptor_write_waitrequest
	wire  [31:0] sgdma_rx_descriptor_write_address;                                 // sgdma_rx:descriptor_write_address -> mm_interconnect_0:sgdma_rx_descriptor_write_address
	wire         sgdma_rx_descriptor_write_write;                                   // sgdma_rx:descriptor_write_write -> mm_interconnect_0:sgdma_rx_descriptor_write_write
	wire  [31:0] sgdma_rx_descriptor_write_writedata;                               // sgdma_rx:descriptor_write_writedata -> mm_interconnect_0:sgdma_rx_descriptor_write_writedata
	wire         sgdma_tx_descriptor_write_waitrequest;                             // mm_interconnect_0:sgdma_tx_descriptor_write_waitrequest -> sgdma_tx:descriptor_write_waitrequest
	wire  [31:0] sgdma_tx_descriptor_write_address;                                 // sgdma_tx:descriptor_write_address -> mm_interconnect_0:sgdma_tx_descriptor_write_address
	wire         sgdma_tx_descriptor_write_write;                                   // sgdma_tx:descriptor_write_write -> mm_interconnect_0:sgdma_tx_descriptor_write_write
	wire  [31:0] sgdma_tx_descriptor_write_writedata;                               // sgdma_tx:descriptor_write_writedata -> mm_interconnect_0:sgdma_tx_descriptor_write_writedata
	wire  [31:0] nios2_gen2_instruction_master_readdata;                            // mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	wire         nios2_gen2_instruction_master_waitrequest;                         // mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	wire  [29:0] nios2_gen2_instruction_master_address;                             // nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
	wire         nios2_gen2_instruction_master_read;                                // nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
	wire         nios2_gen2_instruction_master_readdatavalid;                       // mm_interconnect_0:nios2_gen2_instruction_master_readdatavalid -> nios2_gen2:i_readdatavalid
	wire  [31:0] sgdma_tx_m_read_readdata;                                          // mm_interconnect_0:sgdma_tx_m_read_readdata -> sgdma_tx:m_read_readdata
	wire         sgdma_tx_m_read_waitrequest;                                       // mm_interconnect_0:sgdma_tx_m_read_waitrequest -> sgdma_tx:m_read_waitrequest
	wire  [31:0] sgdma_tx_m_read_address;                                           // sgdma_tx:m_read_address -> mm_interconnect_0:sgdma_tx_m_read_address
	wire         sgdma_tx_m_read_read;                                              // sgdma_tx:m_read_read -> mm_interconnect_0:sgdma_tx_m_read_read
	wire         sgdma_tx_m_read_readdatavalid;                                     // mm_interconnect_0:sgdma_tx_m_read_readdatavalid -> sgdma_tx:m_read_readdatavalid
	wire         sgdma_rx_m_write_waitrequest;                                      // mm_interconnect_0:sgdma_rx_m_write_waitrequest -> sgdma_rx:m_write_waitrequest
	wire  [31:0] sgdma_rx_m_write_address;                                          // sgdma_rx:m_write_address -> mm_interconnect_0:sgdma_rx_m_write_address
	wire   [3:0] sgdma_rx_m_write_byteenable;                                       // sgdma_rx:m_write_byteenable -> mm_interconnect_0:sgdma_rx_m_write_byteenable
	wire         sgdma_rx_m_write_write;                                            // sgdma_rx:m_write_write -> mm_interconnect_0:sgdma_rx_m_write_write
	wire  [31:0] sgdma_rx_m_write_writedata;                                        // sgdma_rx:m_write_writedata -> mm_interconnect_0:sgdma_rx_m_write_writedata
	wire  [31:0] mm_interconnect_0_tse_mac_control_port_readdata;                   // tse_mac:reg_data_out -> mm_interconnect_0:tse_mac_control_port_readdata
	wire         mm_interconnect_0_tse_mac_control_port_waitrequest;                // tse_mac:reg_busy -> mm_interconnect_0:tse_mac_control_port_waitrequest
	wire   [7:0] mm_interconnect_0_tse_mac_control_port_address;                    // mm_interconnect_0:tse_mac_control_port_address -> tse_mac:reg_addr
	wire         mm_interconnect_0_tse_mac_control_port_read;                       // mm_interconnect_0:tse_mac_control_port_read -> tse_mac:reg_rd
	wire         mm_interconnect_0_tse_mac_control_port_write;                      // mm_interconnect_0:tse_mac_control_port_write -> tse_mac:reg_wr
	wire  [31:0] mm_interconnect_0_tse_mac_control_port_writedata;                  // mm_interconnect_0:tse_mac_control_port_writedata -> tse_mac:reg_data_in
	wire         mm_interconnect_0_sgdma_tx_csr_chipselect;                         // mm_interconnect_0:sgdma_tx_csr_chipselect -> sgdma_tx:csr_chipselect
	wire  [31:0] mm_interconnect_0_sgdma_tx_csr_readdata;                           // sgdma_tx:csr_readdata -> mm_interconnect_0:sgdma_tx_csr_readdata
	wire   [3:0] mm_interconnect_0_sgdma_tx_csr_address;                            // mm_interconnect_0:sgdma_tx_csr_address -> sgdma_tx:csr_address
	wire         mm_interconnect_0_sgdma_tx_csr_read;                               // mm_interconnect_0:sgdma_tx_csr_read -> sgdma_tx:csr_read
	wire         mm_interconnect_0_sgdma_tx_csr_write;                              // mm_interconnect_0:sgdma_tx_csr_write -> sgdma_tx:csr_write
	wire  [31:0] mm_interconnect_0_sgdma_tx_csr_writedata;                          // mm_interconnect_0:sgdma_tx_csr_writedata -> sgdma_tx:csr_writedata
	wire         mm_interconnect_0_sgdma_rx_csr_chipselect;                         // mm_interconnect_0:sgdma_rx_csr_chipselect -> sgdma_rx:csr_chipselect
	wire  [31:0] mm_interconnect_0_sgdma_rx_csr_readdata;                           // sgdma_rx:csr_readdata -> mm_interconnect_0:sgdma_rx_csr_readdata
	wire   [3:0] mm_interconnect_0_sgdma_rx_csr_address;                            // mm_interconnect_0:sgdma_rx_csr_address -> sgdma_rx:csr_address
	wire         mm_interconnect_0_sgdma_rx_csr_read;                               // mm_interconnect_0:sgdma_rx_csr_read -> sgdma_rx:csr_read
	wire         mm_interconnect_0_sgdma_rx_csr_write;                              // mm_interconnect_0:sgdma_rx_csr_write -> sgdma_rx:csr_write
	wire  [31:0] mm_interconnect_0_sgdma_rx_csr_writedata;                          // mm_interconnect_0:sgdma_rx_csr_writedata -> sgdma_rx:csr_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata;             // nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest;          // nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess;          // mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_address;              // mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_read;                 // mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable;           // mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_debug_mem_slave_write;                // mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata;            // mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                          // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                           // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_read;                              // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire         mm_interconnect_0_pll_pll_slave_write;                             // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                         // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire  [31:0] mm_interconnect_0_slow_periph_bridge_s0_readdata;                  // slow_periph_bridge:s0_readdata -> mm_interconnect_0:slow_periph_bridge_s0_readdata
	wire         mm_interconnect_0_slow_periph_bridge_s0_waitrequest;               // slow_periph_bridge:s0_waitrequest -> mm_interconnect_0:slow_periph_bridge_s0_waitrequest
	wire         mm_interconnect_0_slow_periph_bridge_s0_debugaccess;               // mm_interconnect_0:slow_periph_bridge_s0_debugaccess -> slow_periph_bridge:s0_debugaccess
	wire   [9:0] mm_interconnect_0_slow_periph_bridge_s0_address;                   // mm_interconnect_0:slow_periph_bridge_s0_address -> slow_periph_bridge:s0_address
	wire         mm_interconnect_0_slow_periph_bridge_s0_read;                      // mm_interconnect_0:slow_periph_bridge_s0_read -> slow_periph_bridge:s0_read
	wire   [3:0] mm_interconnect_0_slow_periph_bridge_s0_byteenable;                // mm_interconnect_0:slow_periph_bridge_s0_byteenable -> slow_periph_bridge:s0_byteenable
	wire         mm_interconnect_0_slow_periph_bridge_s0_readdatavalid;             // slow_periph_bridge:s0_readdatavalid -> mm_interconnect_0:slow_periph_bridge_s0_readdatavalid
	wire         mm_interconnect_0_slow_periph_bridge_s0_write;                     // mm_interconnect_0:slow_periph_bridge_s0_write -> slow_periph_bridge:s0_write
	wire  [31:0] mm_interconnect_0_slow_periph_bridge_s0_writedata;                 // mm_interconnect_0:slow_periph_bridge_s0_writedata -> slow_periph_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_slow_periph_bridge_s0_burstcount;                // mm_interconnect_0:slow_periph_bridge_s0_burstcount -> slow_periph_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata;          // mm_clock_crossing_bridge_0:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_readdata
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest;       // mm_clock_crossing_bridge_0:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_waitrequest
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess;       // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_debugaccess -> mm_clock_crossing_bridge_0:s0_debugaccess
	wire  [28:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address;           // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_address -> mm_clock_crossing_bridge_0:s0_address
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read;              // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_read -> mm_clock_crossing_bridge_0:s0_read
	wire   [3:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable;        // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_byteenable -> mm_clock_crossing_bridge_0:s0_byteenable
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid;     // mm_clock_crossing_bridge_0:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_0_s0_readdatavalid
	wire         mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write;             // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_write -> mm_clock_crossing_bridge_0:s0_write
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata;         // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_writedata -> mm_clock_crossing_bridge_0:s0_writedata
	wire   [0:0] mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount;        // mm_interconnect_0:mm_clock_crossing_bridge_0_s0_burstcount -> mm_clock_crossing_bridge_0:s0_burstcount
	wire         mm_interconnect_0_descriptor_memory_s1_chipselect;                 // mm_interconnect_0:descriptor_memory_s1_chipselect -> descriptor_memory:chipselect
	wire  [31:0] mm_interconnect_0_descriptor_memory_s1_readdata;                   // descriptor_memory:readdata -> mm_interconnect_0:descriptor_memory_s1_readdata
	wire   [9:0] mm_interconnect_0_descriptor_memory_s1_address;                    // mm_interconnect_0:descriptor_memory_s1_address -> descriptor_memory:address
	wire   [3:0] mm_interconnect_0_descriptor_memory_s1_byteenable;                 // mm_interconnect_0:descriptor_memory_s1_byteenable -> descriptor_memory:byteenable
	wire         mm_interconnect_0_descriptor_memory_s1_write;                      // mm_interconnect_0:descriptor_memory_s1_write -> descriptor_memory:write
	wire  [31:0] mm_interconnect_0_descriptor_memory_s1_writedata;                  // mm_interconnect_0:descriptor_memory_s1_writedata -> descriptor_memory:writedata
	wire         mm_interconnect_0_descriptor_memory_s1_clken;                      // mm_interconnect_0:descriptor_memory_s1_clken -> descriptor_memory:clken
	wire         slow_periph_bridge_m0_waitrequest;                                 // mm_interconnect_1:slow_periph_bridge_m0_waitrequest -> slow_periph_bridge:m0_waitrequest
	wire  [31:0] slow_periph_bridge_m0_readdata;                                    // mm_interconnect_1:slow_periph_bridge_m0_readdata -> slow_periph_bridge:m0_readdata
	wire         slow_periph_bridge_m0_debugaccess;                                 // slow_periph_bridge:m0_debugaccess -> mm_interconnect_1:slow_periph_bridge_m0_debugaccess
	wire   [9:0] slow_periph_bridge_m0_address;                                     // slow_periph_bridge:m0_address -> mm_interconnect_1:slow_periph_bridge_m0_address
	wire         slow_periph_bridge_m0_read;                                        // slow_periph_bridge:m0_read -> mm_interconnect_1:slow_periph_bridge_m0_read
	wire   [3:0] slow_periph_bridge_m0_byteenable;                                  // slow_periph_bridge:m0_byteenable -> mm_interconnect_1:slow_periph_bridge_m0_byteenable
	wire         slow_periph_bridge_m0_readdatavalid;                               // mm_interconnect_1:slow_periph_bridge_m0_readdatavalid -> slow_periph_bridge:m0_readdatavalid
	wire  [31:0] slow_periph_bridge_m0_writedata;                                   // slow_periph_bridge:m0_writedata -> mm_interconnect_1:slow_periph_bridge_m0_writedata
	wire         slow_periph_bridge_m0_write;                                       // slow_periph_bridge:m0_write -> mm_interconnect_1:slow_periph_bridge_m0_write
	wire   [0:0] slow_periph_bridge_m0_burstcount;                                  // slow_periph_bridge:m0_burstcount -> mm_interconnect_1:slow_periph_bridge_m0_burstcount
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect;          // mm_interconnect_1:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata;            // jtag_uart:av_readdata -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest;         // jtag_uart:av_waitrequest -> mm_interconnect_1:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_address;             // mm_interconnect_1:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_read;                // mm_interconnect_1:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_1_jtag_uart_avalon_jtag_slave_write;               // mm_interconnect_1:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata;           // mm_interconnect_1:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_1_performance_counter_control_slave_readdata;      // performance_counter:readdata -> mm_interconnect_1:performance_counter_control_slave_readdata
	wire   [3:0] mm_interconnect_1_performance_counter_control_slave_address;       // mm_interconnect_1:performance_counter_control_slave_address -> performance_counter:address
	wire         mm_interconnect_1_performance_counter_control_slave_begintransfer; // mm_interconnect_1:performance_counter_control_slave_begintransfer -> performance_counter:begintransfer
	wire         mm_interconnect_1_performance_counter_control_slave_write;         // mm_interconnect_1:performance_counter_control_slave_write -> performance_counter:write
	wire  [31:0] mm_interconnect_1_performance_counter_control_slave_writedata;     // mm_interconnect_1:performance_counter_control_slave_writedata -> performance_counter:writedata
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;                    // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;                     // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_1_sys_timer_s1_chipselect;                         // mm_interconnect_1:sys_timer_s1_chipselect -> sys_timer:chipselect
	wire  [15:0] mm_interconnect_1_sys_timer_s1_readdata;                           // sys_timer:readdata -> mm_interconnect_1:sys_timer_s1_readdata
	wire   [2:0] mm_interconnect_1_sys_timer_s1_address;                            // mm_interconnect_1:sys_timer_s1_address -> sys_timer:address
	wire         mm_interconnect_1_sys_timer_s1_write;                              // mm_interconnect_1:sys_timer_s1_write -> sys_timer:write_n
	wire  [15:0] mm_interconnect_1_sys_timer_s1_writedata;                          // mm_interconnect_1:sys_timer_s1_writedata -> sys_timer:writedata
	wire         mm_interconnect_1_high_res_timer_s1_chipselect;                    // mm_interconnect_1:high_res_timer_s1_chipselect -> high_res_timer:chipselect
	wire  [15:0] mm_interconnect_1_high_res_timer_s1_readdata;                      // high_res_timer:readdata -> mm_interconnect_1:high_res_timer_s1_readdata
	wire   [2:0] mm_interconnect_1_high_res_timer_s1_address;                       // mm_interconnect_1:high_res_timer_s1_address -> high_res_timer:address
	wire         mm_interconnect_1_high_res_timer_s1_write;                         // mm_interconnect_1:high_res_timer_s1_write -> high_res_timer:write_n
	wire  [15:0] mm_interconnect_1_high_res_timer_s1_writedata;                     // mm_interconnect_1:high_res_timer_s1_writedata -> high_res_timer:writedata
	wire         mm_interconnect_1_led_pio_s1_chipselect;                           // mm_interconnect_1:led_pio_s1_chipselect -> led_pio:chipselect
	wire  [31:0] mm_interconnect_1_led_pio_s1_readdata;                             // led_pio:readdata -> mm_interconnect_1:led_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_led_pio_s1_address;                              // mm_interconnect_1:led_pio_s1_address -> led_pio:address
	wire         mm_interconnect_1_led_pio_s1_write;                                // mm_interconnect_1:led_pio_s1_write -> led_pio:write_n
	wire  [31:0] mm_interconnect_1_led_pio_s1_writedata;                            // mm_interconnect_1:led_pio_s1_writedata -> led_pio:writedata
	wire         mm_interconnect_1_dipsw_pio_s1_chipselect;                         // mm_interconnect_1:dipsw_pio_s1_chipselect -> dipsw_pio:chipselect
	wire  [31:0] mm_interconnect_1_dipsw_pio_s1_readdata;                           // dipsw_pio:readdata -> mm_interconnect_1:dipsw_pio_s1_readdata
	wire   [1:0] mm_interconnect_1_dipsw_pio_s1_address;                            // mm_interconnect_1:dipsw_pio_s1_address -> dipsw_pio:address
	wire         mm_interconnect_1_dipsw_pio_s1_write;                              // mm_interconnect_1:dipsw_pio_s1_write -> dipsw_pio:write_n
	wire  [31:0] mm_interconnect_1_dipsw_pio_s1_writedata;                          // mm_interconnect_1:dipsw_pio_s1_writedata -> dipsw_pio:writedata
	wire  [31:0] mm_interconnect_1_user_pio_pushbtn_s1_readdata;                    // user_pio_pushbtn:readdata -> mm_interconnect_1:user_pio_pushbtn_s1_readdata
	wire   [1:0] mm_interconnect_1_user_pio_pushbtn_s1_address;                     // mm_interconnect_1:user_pio_pushbtn_s1_address -> user_pio_pushbtn:address
	wire         mm_interconnect_1_nenet_reg_reset_s1_chipselect;                   // mm_interconnect_1:nENET_reg_reset_s1_chipselect -> nENET_reg_reset:chipselect
	wire  [31:0] mm_interconnect_1_nenet_reg_reset_s1_readdata;                     // nENET_reg_reset:readdata -> mm_interconnect_1:nENET_reg_reset_s1_readdata
	wire   [1:0] mm_interconnect_1_nenet_reg_reset_s1_address;                      // mm_interconnect_1:nENET_reg_reset_s1_address -> nENET_reg_reset:address
	wire         mm_interconnect_1_nenet_reg_reset_s1_write;                        // mm_interconnect_1:nENET_reg_reset_s1_write -> nENET_reg_reset:write_n
	wire  [31:0] mm_interconnect_1_nenet_reg_reset_s1_writedata;                    // mm_interconnect_1:nENET_reg_reset_s1_writedata -> nENET_reg_reset:writedata
	wire  [31:0] mm_interconnect_1_ddr3_status_s1_readdata;                         // ddr3_status:readdata -> mm_interconnect_1:ddr3_status_s1_readdata
	wire   [1:0] mm_interconnect_1_ddr3_status_s1_address;                          // mm_interconnect_1:ddr3_status_s1_address -> ddr3_status:address
	wire         mm_clock_crossing_bridge_0_m0_waitrequest;                         // mm_interconnect_2:mm_clock_crossing_bridge_0_m0_waitrequest -> mm_clock_crossing_bridge_0:m0_waitrequest
	wire  [31:0] mm_clock_crossing_bridge_0_m0_readdata;                            // mm_interconnect_2:mm_clock_crossing_bridge_0_m0_readdata -> mm_clock_crossing_bridge_0:m0_readdata
	wire         mm_clock_crossing_bridge_0_m0_debugaccess;                         // mm_clock_crossing_bridge_0:m0_debugaccess -> mm_interconnect_2:mm_clock_crossing_bridge_0_m0_debugaccess
	wire  [28:0] mm_clock_crossing_bridge_0_m0_address;                             // mm_clock_crossing_bridge_0:m0_address -> mm_interconnect_2:mm_clock_crossing_bridge_0_m0_address
	wire         mm_clock_crossing_bridge_0_m0_read;                                // mm_clock_crossing_bridge_0:m0_read -> mm_interconnect_2:mm_clock_crossing_bridge_0_m0_read
	wire   [3:0] mm_clock_crossing_bridge_0_m0_byteenable;                          // mm_clock_crossing_bridge_0:m0_byteenable -> mm_interconnect_2:mm_clock_crossing_bridge_0_m0_byteenable
	wire         mm_clock_crossing_bridge_0_m0_readdatavalid;                       // mm_interconnect_2:mm_clock_crossing_bridge_0_m0_readdatavalid -> mm_clock_crossing_bridge_0:m0_readdatavalid
	wire  [31:0] mm_clock_crossing_bridge_0_m0_writedata;                           // mm_clock_crossing_bridge_0:m0_writedata -> mm_interconnect_2:mm_clock_crossing_bridge_0_m0_writedata
	wire         mm_clock_crossing_bridge_0_m0_write;                               // mm_clock_crossing_bridge_0:m0_write -> mm_interconnect_2:mm_clock_crossing_bridge_0_m0_write
	wire   [0:0] mm_clock_crossing_bridge_0_m0_burstcount;                          // mm_clock_crossing_bridge_0:m0_burstcount -> mm_interconnect_2:mm_clock_crossing_bridge_0_m0_burstcount
	wire         mm_interconnect_2_mem_if_ddr3_emif_avl_beginbursttransfer;         // mm_interconnect_2:mem_if_ddr3_emif_avl_beginbursttransfer -> mem_if_ddr3_emif:avl_burstbegin
	wire  [63:0] mm_interconnect_2_mem_if_ddr3_emif_avl_readdata;                   // mem_if_ddr3_emif:avl_rdata -> mm_interconnect_2:mem_if_ddr3_emif_avl_readdata
	wire         mm_interconnect_2_mem_if_ddr3_emif_avl_waitrequest;                // mem_if_ddr3_emif:avl_ready -> mm_interconnect_2:mem_if_ddr3_emif_avl_waitrequest
	wire  [25:0] mm_interconnect_2_mem_if_ddr3_emif_avl_address;                    // mm_interconnect_2:mem_if_ddr3_emif_avl_address -> mem_if_ddr3_emif:avl_addr
	wire         mm_interconnect_2_mem_if_ddr3_emif_avl_read;                       // mm_interconnect_2:mem_if_ddr3_emif_avl_read -> mem_if_ddr3_emif:avl_read_req
	wire   [7:0] mm_interconnect_2_mem_if_ddr3_emif_avl_byteenable;                 // mm_interconnect_2:mem_if_ddr3_emif_avl_byteenable -> mem_if_ddr3_emif:avl_be
	wire         mm_interconnect_2_mem_if_ddr3_emif_avl_readdatavalid;              // mem_if_ddr3_emif:avl_rdata_valid -> mm_interconnect_2:mem_if_ddr3_emif_avl_readdatavalid
	wire         mm_interconnect_2_mem_if_ddr3_emif_avl_write;                      // mm_interconnect_2:mem_if_ddr3_emif_avl_write -> mem_if_ddr3_emif:avl_write_req
	wire  [63:0] mm_interconnect_2_mem_if_ddr3_emif_avl_writedata;                  // mm_interconnect_2:mem_if_ddr3_emif_avl_writedata -> mem_if_ddr3_emif:avl_wdata
	wire   [2:0] mm_interconnect_2_mem_if_ddr3_emif_avl_burstcount;                 // mm_interconnect_2:mem_if_ddr3_emif_avl_burstcount -> mem_if_ddr3_emif:avl_size
	wire         irq_mapper_receiver0_irq;                                          // sgdma_tx:csr_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                          // sgdma_rx:csr_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver4_irq;                                          // jtag_uart:av_irq -> irq_mapper:receiver4_irq
	wire  [31:0] nios2_gen2_irq_irq;                                                // irq_mapper:sender_irq -> nios2_gen2:irq
	wire         irq_mapper_receiver2_irq;                                          // irq_synchronizer:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                     // sys_timer:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver3_irq;                                          // irq_synchronizer_001:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                 // high_res_timer:irq -> irq_synchronizer_001:receiver_irq
	wire         tse_mac_receive_valid;                                             // tse_mac:ff_rx_dval -> avalon_st_adapter:in_0_valid
	wire  [31:0] tse_mac_receive_data;                                              // tse_mac:ff_rx_data -> avalon_st_adapter:in_0_data
	wire         tse_mac_receive_ready;                                             // avalon_st_adapter:in_0_ready -> tse_mac:ff_rx_rdy
	wire         tse_mac_receive_startofpacket;                                     // tse_mac:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	wire         tse_mac_receive_endofpacket;                                       // tse_mac:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	wire   [5:0] tse_mac_receive_error;                                             // tse_mac:rx_err -> avalon_st_adapter:in_0_error
	wire   [1:0] tse_mac_receive_empty;                                             // tse_mac:ff_rx_mod -> avalon_st_adapter:in_0_empty
	wire         avalon_st_adapter_out_0_valid;                                     // avalon_st_adapter:out_0_valid -> sgdma_rx:in_valid
	wire  [31:0] avalon_st_adapter_out_0_data;                                      // avalon_st_adapter:out_0_data -> sgdma_rx:in_data
	wire         avalon_st_adapter_out_0_ready;                                     // sgdma_rx:in_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                             // avalon_st_adapter:out_0_startofpacket -> sgdma_rx:in_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                               // avalon_st_adapter:out_0_endofpacket -> sgdma_rx:in_endofpacket
	wire   [5:0] avalon_st_adapter_out_0_error;                                     // avalon_st_adapter:out_0_error -> sgdma_rx:in_error
	wire   [1:0] avalon_st_adapter_out_0_empty;                                     // avalon_st_adapter:out_0_empty -> sgdma_rx:in_empty
	wire         rst_controller_reset_out_reset;                                    // rst_controller:reset_out -> [ddr3_status:reset_n, dipsw_pio:reset_n, high_res_timer:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, led_pio:reset_n, mm_interconnect_1:slow_periph_bridge_m0_reset_reset_bridge_in_reset_reset, nENET_reg_reset:reset_n, performance_counter:reset_n, slow_periph_bridge:m0_reset, sys_timer:reset_n, sysid:reset_n, user_pio_pushbtn:reset_n]
	wire         rst_controller_001_reset_out_reset;                                // rst_controller_001:reset_out -> [avalon_st_adapter:in_rst_0_reset, descriptor_memory:reset, mm_interconnect_0:sgdma_rx_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sgdma_rx:system_reset_n, sgdma_tx:system_reset_n, slow_periph_bridge:s0_reset, tse_mac:reset]
	wire         rst_controller_001_reset_out_reset_req;                            // rst_controller_001:reset_req -> [descriptor_memory:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                                // rst_controller_002:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, jtag_uart:rst_n, mm_clock_crossing_bridge_0:s0_reset, mm_interconnect_0:nios2_gen2_reset_reset_bridge_in_reset_reset, mm_interconnect_1:jtag_uart_reset_reset_bridge_in_reset_reset, nios2_gen2:reset_n, rst_translator_001:in_reset]
	wire         rst_controller_002_reset_out_reset_req;                            // rst_controller_002:reset_req -> [nios2_gen2:reset_req, rst_translator_001:reset_req_in]
	wire         nios2_gen2_debug_reset_request_reset;                              // nios2_gen2:debug_reset_request -> [rst_controller_002:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in1, rst_controller_005:reset_in1]
	wire         rst_controller_003_reset_out_reset;                                // rst_controller_003:reset_out -> mem_if_ddr3_emif:global_reset_n
	wire         rst_controller_004_reset_out_reset;                                // rst_controller_004:reset_out -> mem_if_ddr3_emif:soft_reset_n
	wire         rst_controller_005_reset_out_reset;                                // rst_controller_005:reset_out -> [mm_clock_crossing_bridge_0:m0_reset, mm_interconnect_2:mem_if_ddr3_emif_soft_reset_reset_bridge_in_reset_reset, mm_interconnect_2:mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_006_reset_out_reset;                                // rst_controller_006:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]

	DECA_Qsys_ddr3_status ddr3_status (
		.clk      (pll_c2_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_1_ddr3_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_ddr3_status_s1_readdata), //                    .readdata
		.in_port  (ddr3_status_external_connection_export)     // external_connection.export
	);

	DECA_Qsys_descriptor_memory descriptor_memory (
		.clk        (pll_c0_clk),                                        //   clk1.clk
		.address    (mm_interconnect_0_descriptor_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_descriptor_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_descriptor_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_descriptor_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_descriptor_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_descriptor_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_descriptor_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req)             //       .reset_req
	);

	DECA_Qsys_dipsw_pio dipsw_pio (
		.clk        (pll_c2_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_1_dipsw_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_dipsw_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_dipsw_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_dipsw_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_dipsw_pio_s1_readdata),   //                    .readdata
		.in_port    (dipsw_pio_export)                           // external_connection.export
	);

	DECA_Qsys_high_res_timer high_res_timer (
		.clk        (pll_c2_clk),                                     //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                // reset.reset_n
		.address    (mm_interconnect_1_high_res_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_high_res_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_high_res_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_high_res_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_high_res_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)               //   irq.irq
	);

	DECA_Qsys_jtag_uart jtag_uart (
		.clk            (pll_c0_clk),                                                //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver4_irq)                                   //               irq.irq
	);

	DECA_Qsys_led_pio led_pio (
		.clk        (pll_c2_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_led_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_led_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_led_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_led_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_led_pio_s1_readdata),   //                    .readdata
		.out_port   (led_pio_export)                           // external_connection.export
	);

	DECA_Qsys_mem_if_ddr3_emif mem_if_ddr3_emif (
		.pll_ref_clk        (mem_if_ddr3_emif_pll_ref_clk_clk),                          //      pll_ref_clk.clk
		.global_reset_n     (~rst_controller_003_reset_out_reset),                       //     global_reset.reset_n
		.soft_reset_n       (~rst_controller_004_reset_out_reset),                       //       soft_reset.reset_n
		.afi_clk            (mem_if_ddr3_emif_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk       (),                                                          //     afi_half_clk.clk
		.afi_reset_n        (),                                                          //        afi_reset.reset_n
		.afi_reset_export_n (),                                                          // afi_reset_export.reset_n
		.mem_a              (memory_mem_a),                                              //           memory.mem_a
		.mem_ba             (memory_mem_ba),                                             //                 .mem_ba
		.mem_ck             (memory_mem_ck),                                             //                 .mem_ck
		.mem_ck_n           (memory_mem_ck_n),                                           //                 .mem_ck_n
		.mem_cke            (memory_mem_cke),                                            //                 .mem_cke
		.mem_cs_n           (memory_mem_cs_n),                                           //                 .mem_cs_n
		.mem_dm             (memory_mem_dm),                                             //                 .mem_dm
		.mem_ras_n          (memory_mem_ras_n),                                          //                 .mem_ras_n
		.mem_cas_n          (memory_mem_cas_n),                                          //                 .mem_cas_n
		.mem_we_n           (memory_mem_we_n),                                           //                 .mem_we_n
		.mem_reset_n        (memory_mem_reset_n),                                        //                 .mem_reset_n
		.mem_dq             (memory_mem_dq),                                             //                 .mem_dq
		.mem_dqs            (memory_mem_dqs),                                            //                 .mem_dqs
		.mem_dqs_n          (memory_mem_dqs_n),                                          //                 .mem_dqs_n
		.mem_odt            (memory_mem_odt),                                            //                 .mem_odt
		.avl_ready          (mm_interconnect_2_mem_if_ddr3_emif_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin     (mm_interconnect_2_mem_if_ddr3_emif_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr           (mm_interconnect_2_mem_if_ddr3_emif_avl_address),            //                 .address
		.avl_rdata_valid    (mm_interconnect_2_mem_if_ddr3_emif_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata          (mm_interconnect_2_mem_if_ddr3_emif_avl_readdata),           //                 .readdata
		.avl_wdata          (mm_interconnect_2_mem_if_ddr3_emif_avl_writedata),          //                 .writedata
		.avl_be             (mm_interconnect_2_mem_if_ddr3_emif_avl_byteenable),         //                 .byteenable
		.avl_read_req       (mm_interconnect_2_mem_if_ddr3_emif_avl_read),               //                 .read
		.avl_write_req      (mm_interconnect_2_mem_if_ddr3_emif_avl_write),              //                 .write
		.avl_size           (mm_interconnect_2_mem_if_ddr3_emif_avl_burstcount),         //                 .burstcount
		.local_init_done    (mem_if_ddr3_emif_status_local_init_done),                   //           status.local_init_done
		.local_cal_success  (mem_if_ddr3_emif_status_local_cal_success),                 //                 .local_cal_success
		.local_cal_fail     (mem_if_ddr3_emif_status_local_cal_fail),                    //                 .local_cal_fail
		.pll_mem_clk        (mem_if_ddr3_emif_pll_sharing_pll_mem_clk),                  //      pll_sharing.pll_mem_clk
		.pll_write_clk      (mem_if_ddr3_emif_pll_sharing_pll_write_clk),                //                 .pll_write_clk
		.pll_locked         (mem_if_ddr3_emif_pll_sharing_pll_locked),                   //                 .pll_locked
		.pll_capture0_clk   (mem_if_ddr3_emif_pll_sharing_pll_capture0_clk),             //                 .pll_capture0_clk
		.pll_capture1_clk   (mem_if_ddr3_emif_pll_sharing_pll_capture1_clk)              //                 .pll_capture1_clk
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (29),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (16),
		.RESPONSE_FIFO_DEPTH (16),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge_0 (
		.m0_clk           (mem_if_ddr3_emif_afi_clk_clk),                                  //   m0_clk.clk
		.m0_reset         (rst_controller_005_reset_out_reset),                            // m0_reset.reset
		.s0_clk           (pll_c0_clk),                                                    //   s0_clk.clk
		.s0_reset         (rst_controller_002_reset_out_reset),                            // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_0_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_0_m0_readdata),                        //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_0_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_0_m0_burstcount),                      //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_0_m0_writedata),                       //         .writedata
		.m0_address       (mm_clock_crossing_bridge_0_m0_address),                         //         .address
		.m0_write         (mm_clock_crossing_bridge_0_m0_write),                           //         .write
		.m0_read          (mm_clock_crossing_bridge_0_m0_read),                            //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_0_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_0_m0_debugaccess)                      //         .debugaccess
	);

	DECA_Qsys_nENET_reg_reset nenet_reg_reset (
		.clk        (pll_c2_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_1_nenet_reg_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_nenet_reg_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_nenet_reg_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_nenet_reg_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_nenet_reg_reset_s1_readdata),   //                    .readdata
		.out_port   (nenet_reg_reset_export)                           // external_connection.export
	);

	DECA_Qsys_nios2_gen2 nios2_gen2 (
		.clk                                 (pll_c0_clk),                                               //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_gen2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	DECA_Qsys_performance_counter performance_counter (
		.clk           (pll_c2_clk),                                                        //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                   //         reset.reset_n
		.address       (mm_interconnect_1_performance_counter_control_slave_address),       // control_slave.address
		.begintransfer (mm_interconnect_1_performance_counter_control_slave_begintransfer), //              .begintransfer
		.readdata      (mm_interconnect_1_performance_counter_control_slave_readdata),      //              .readdata
		.write         (mm_interconnect_1_performance_counter_control_slave_write),         //              .write
		.writedata     (mm_interconnect_1_performance_counter_control_slave_writedata)      //              .writedata
	);

	DECA_Qsys_pll pll (
		.clk       (clk_clk),                                   //       inclk_interface.clk
		.reset     (rst_controller_006_reset_out_reset),        // inclk_interface_reset.reset
		.read      (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0        (pll_c0_clk),                                //                    c0.clk
		.c1        (),                                          //                    c1.clk
		.c2        (pll_c2_clk),                                //                    c2.clk
		.c3        (),                                          //                    c3.clk
		.areset    (pll_areset_conduit_export),                 //        areset_conduit.export
		.locked    (pll_locked_conduit_export),                 //        locked_conduit.export
		.phasedone (pll_phasedone_conduit_export)               //     phasedone_conduit.export
	);

	DECA_Qsys_sgdma_rx sgdma_rx (
		.clk                           (pll_c0_clk),                                //              clk.clk
		.system_reset_n                (~rst_controller_001_reset_out_reset),       //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_rx_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_rx_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_rx_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_rx_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_rx_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_rx_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_rx_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_rx_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_rx_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_rx_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_rx_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_rx_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_rx_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_rx_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_rx_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver1_irq),                  //          csr_irq.irq
		.in_startofpacket              (avalon_st_adapter_out_0_startofpacket),     //               in.startofpacket
		.in_endofpacket                (avalon_st_adapter_out_0_endofpacket),       //                 .endofpacket
		.in_data                       (avalon_st_adapter_out_0_data),              //                 .data
		.in_valid                      (avalon_st_adapter_out_0_valid),             //                 .valid
		.in_ready                      (avalon_st_adapter_out_0_ready),             //                 .ready
		.in_empty                      (avalon_st_adapter_out_0_empty),             //                 .empty
		.in_error                      (avalon_st_adapter_out_0_error),             //                 .error
		.m_write_waitrequest           (sgdma_rx_m_write_waitrequest),              //          m_write.waitrequest
		.m_write_address               (sgdma_rx_m_write_address),                  //                 .address
		.m_write_write                 (sgdma_rx_m_write_write),                    //                 .write
		.m_write_writedata             (sgdma_rx_m_write_writedata),                //                 .writedata
		.m_write_byteenable            (sgdma_rx_m_write_byteenable)                //                 .byteenable
	);

	DECA_Qsys_sgdma_tx sgdma_tx (
		.clk                           (pll_c0_clk),                                //              clk.clk
		.system_reset_n                (~rst_controller_001_reset_out_reset),       //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_tx_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_tx_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_tx_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_tx_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_tx_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_tx_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_tx_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_tx_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_tx_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_tx_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_tx_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_tx_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_tx_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_tx_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_tx_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),                  //          csr_irq.irq
		.m_read_readdata               (sgdma_tx_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (sgdma_tx_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (sgdma_tx_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (sgdma_tx_m_read_address),                   //                 .address
		.m_read_read                   (sgdma_tx_m_read_read),                      //                 .read
		.out_data                      (sgdma_tx_out_data),                         //              out.data
		.out_valid                     (sgdma_tx_out_valid),                        //                 .valid
		.out_ready                     (sgdma_tx_out_ready),                        //                 .ready
		.out_endofpacket               (sgdma_tx_out_endofpacket),                  //                 .endofpacket
		.out_startofpacket             (sgdma_tx_out_startofpacket),                //                 .startofpacket
		.out_empty                     (sgdma_tx_out_empty),                        //                 .empty
		.out_error                     (sgdma_tx_out_error)                         //                 .error
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) slow_periph_bridge (
		.m0_clk           (pll_c2_clk),                                            //   m0_clk.clk
		.m0_reset         (rst_controller_reset_out_reset),                        // m0_reset.reset
		.s0_clk           (pll_c0_clk),                                            //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                    // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_slow_periph_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_slow_periph_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_slow_periph_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_slow_periph_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_slow_periph_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_slow_periph_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_slow_periph_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_slow_periph_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_slow_periph_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_slow_periph_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (slow_periph_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (slow_periph_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (slow_periph_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (slow_periph_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (slow_periph_bridge_m0_writedata),                       //         .writedata
		.m0_address       (slow_periph_bridge_m0_address),                         //         .address
		.m0_write         (slow_periph_bridge_m0_write),                           //         .write
		.m0_read          (slow_periph_bridge_m0_read),                            //         .read
		.m0_byteenable    (slow_periph_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (slow_periph_bridge_m0_debugaccess)                      //         .debugaccess
	);

	DECA_Qsys_sys_timer sys_timer (
		.clk        (pll_c2_clk),                                //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_1_sys_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_sys_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_sys_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_sys_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_sys_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)              //   irq.irq
	);

	DECA_Qsys_sysid sysid (
		.clock    (pll_c2_clk),                                     //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	DECA_Qsys_tse_mac tse_mac (
		.clk           (pll_c0_clk),                                         // control_port_clock_connection.clk
		.reset         (rst_controller_001_reset_out_reset),                 //              reset_connection.reset
		.reg_addr      (mm_interconnect_0_tse_mac_control_port_address),     //                  control_port.address
		.reg_data_out  (mm_interconnect_0_tse_mac_control_port_readdata),    //                              .readdata
		.reg_rd        (mm_interconnect_0_tse_mac_control_port_read),        //                              .read
		.reg_data_in   (mm_interconnect_0_tse_mac_control_port_writedata),   //                              .writedata
		.reg_wr        (mm_interconnect_0_tse_mac_control_port_write),       //                              .write
		.reg_busy      (mm_interconnect_0_tse_mac_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (tse_mac_pcs_mac_tx_clock_connection_clk),            //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (tse_mac_pcs_mac_rx_clock_connection_clk),            //   pcs_mac_rx_clock_connection.clk
		.set_10        (tse_mac_mac_status_connection_set_10),               //         mac_status_connection.set_10
		.set_1000      (tse_mac_mac_status_connection_set_1000),             //                              .set_1000
		.eth_mode      (tse_mac_mac_status_connection_eth_mode),             //                              .eth_mode
		.ena_10        (tse_mac_mac_status_connection_ena_10),               //                              .ena_10
		.m_rx_d        (tse_mac_mac_mii_connection_mii_rx_d),                //            mac_mii_connection.mii_rx_d
		.m_rx_en       (tse_mac_mac_mii_connection_mii_rx_dv),               //                              .mii_rx_dv
		.m_rx_err      (tse_mac_mac_mii_connection_mii_rx_err),              //                              .mii_rx_err
		.m_tx_d        (tse_mac_mac_mii_connection_mii_tx_d),                //                              .mii_tx_d
		.m_tx_en       (tse_mac_mac_mii_connection_mii_tx_en),               //                              .mii_tx_en
		.m_tx_err      (tse_mac_mac_mii_connection_mii_tx_err),              //                              .mii_tx_err
		.m_rx_crs      (tse_mac_mac_mii_connection_mii_crs),                 //                              .mii_crs
		.m_rx_col      (tse_mac_mac_mii_connection_mii_col),                 //                              .mii_col
		.ff_rx_clk     (pll_c0_clk),                                         //      receive_clock_connection.clk
		.ff_tx_clk     (pll_c0_clk),                                         //     transmit_clock_connection.clk
		.ff_rx_data    (tse_mac_receive_data),                               //                       receive.data
		.ff_rx_eop     (tse_mac_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (tse_mac_receive_error),                              //                              .error
		.ff_rx_mod     (tse_mac_receive_empty),                              //                              .empty
		.ff_rx_rdy     (tse_mac_receive_ready),                              //                              .ready
		.ff_rx_sop     (tse_mac_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (tse_mac_receive_valid),                              //                              .valid
		.ff_tx_data    (sgdma_tx_out_data),                                  //                      transmit.data
		.ff_tx_eop     (sgdma_tx_out_endofpacket),                           //                              .endofpacket
		.ff_tx_err     (sgdma_tx_out_error),                                 //                              .error
		.ff_tx_mod     (sgdma_tx_out_empty),                                 //                              .empty
		.ff_tx_rdy     (sgdma_tx_out_ready),                                 //                              .ready
		.ff_tx_sop     (sgdma_tx_out_startofpacket),                         //                              .startofpacket
		.ff_tx_wren    (sgdma_tx_out_valid),                                 //                              .valid
		.mdc           (tse_mac_mac_mdio_connection_mdc),                    //           mac_mdio_connection.mdc
		.mdio_in       (tse_mac_mac_mdio_connection_mdio_in),                //                              .mdio_in
		.mdio_out      (tse_mac_mac_mdio_connection_mdio_out),               //                              .mdio_out
		.mdio_oen      (tse_mac_mac_mdio_connection_mdio_oen),               //                              .mdio_oen
		.ff_tx_crc_fwd (tse_mac_mac_misc_connection_ff_tx_crc_fwd),          //           mac_misc_connection.ff_tx_crc_fwd
		.ff_tx_septy   (tse_mac_mac_misc_connection_ff_tx_septy),            //                              .ff_tx_septy
		.tx_ff_uflow   (tse_mac_mac_misc_connection_tx_ff_uflow),            //                              .tx_ff_uflow
		.ff_tx_a_full  (tse_mac_mac_misc_connection_ff_tx_a_full),           //                              .ff_tx_a_full
		.ff_tx_a_empty (tse_mac_mac_misc_connection_ff_tx_a_empty),          //                              .ff_tx_a_empty
		.rx_err_stat   (tse_mac_mac_misc_connection_rx_err_stat),            //                              .rx_err_stat
		.rx_frm_type   (tse_mac_mac_misc_connection_rx_frm_type),            //                              .rx_frm_type
		.ff_rx_dsav    (tse_mac_mac_misc_connection_ff_rx_dsav),             //                              .ff_rx_dsav
		.ff_rx_a_full  (tse_mac_mac_misc_connection_ff_rx_a_full),           //                              .ff_rx_a_full
		.ff_rx_a_empty (tse_mac_mac_misc_connection_ff_rx_a_empty)           //                              .ff_rx_a_empty
	);

	DECA_Qsys_user_pio_pushbtn user_pio_pushbtn (
		.clk      (pll_c2_clk),                                     //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address  (mm_interconnect_1_user_pio_pushbtn_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_user_pio_pushbtn_s1_readdata), //                    .readdata
		.in_port  (user_pio_pushbtn_export)                         // external_connection.export
	);

	DECA_Qsys_mm_interconnect_0 mm_interconnect_0 (
		.ext_clk_50_clk_clk                                    (clk_clk),                                                       //                                  ext_clk_50_clk.clk
		.pll_c0_clk                                            (pll_c0_clk),                                                    //                                          pll_c0.clk
		.nios2_gen2_reset_reset_bridge_in_reset_reset          (rst_controller_002_reset_out_reset),                            //          nios2_gen2_reset_reset_bridge_in_reset.reset
		.pll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_006_reset_out_reset),                            // pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.sgdma_rx_reset_reset_bridge_in_reset_reset            (rst_controller_001_reset_out_reset),                            //            sgdma_rx_reset_reset_bridge_in_reset.reset
		.nios2_gen2_data_master_address                        (nios2_gen2_data_master_address),                                //                          nios2_gen2_data_master.address
		.nios2_gen2_data_master_waitrequest                    (nios2_gen2_data_master_waitrequest),                            //                                                .waitrequest
		.nios2_gen2_data_master_byteenable                     (nios2_gen2_data_master_byteenable),                             //                                                .byteenable
		.nios2_gen2_data_master_read                           (nios2_gen2_data_master_read),                                   //                                                .read
		.nios2_gen2_data_master_readdata                       (nios2_gen2_data_master_readdata),                               //                                                .readdata
		.nios2_gen2_data_master_readdatavalid                  (nios2_gen2_data_master_readdatavalid),                          //                                                .readdatavalid
		.nios2_gen2_data_master_write                          (nios2_gen2_data_master_write),                                  //                                                .write
		.nios2_gen2_data_master_writedata                      (nios2_gen2_data_master_writedata),                              //                                                .writedata
		.nios2_gen2_data_master_debugaccess                    (nios2_gen2_data_master_debugaccess),                            //                                                .debugaccess
		.nios2_gen2_instruction_master_address                 (nios2_gen2_instruction_master_address),                         //                   nios2_gen2_instruction_master.address
		.nios2_gen2_instruction_master_waitrequest             (nios2_gen2_instruction_master_waitrequest),                     //                                                .waitrequest
		.nios2_gen2_instruction_master_read                    (nios2_gen2_instruction_master_read),                            //                                                .read
		.nios2_gen2_instruction_master_readdata                (nios2_gen2_instruction_master_readdata),                        //                                                .readdata
		.nios2_gen2_instruction_master_readdatavalid           (nios2_gen2_instruction_master_readdatavalid),                   //                                                .readdatavalid
		.sgdma_rx_descriptor_read_address                      (sgdma_rx_descriptor_read_address),                              //                        sgdma_rx_descriptor_read.address
		.sgdma_rx_descriptor_read_waitrequest                  (sgdma_rx_descriptor_read_waitrequest),                          //                                                .waitrequest
		.sgdma_rx_descriptor_read_read                         (sgdma_rx_descriptor_read_read),                                 //                                                .read
		.sgdma_rx_descriptor_read_readdata                     (sgdma_rx_descriptor_read_readdata),                             //                                                .readdata
		.sgdma_rx_descriptor_read_readdatavalid                (sgdma_rx_descriptor_read_readdatavalid),                        //                                                .readdatavalid
		.sgdma_rx_descriptor_write_address                     (sgdma_rx_descriptor_write_address),                             //                       sgdma_rx_descriptor_write.address
		.sgdma_rx_descriptor_write_waitrequest                 (sgdma_rx_descriptor_write_waitrequest),                         //                                                .waitrequest
		.sgdma_rx_descriptor_write_write                       (sgdma_rx_descriptor_write_write),                               //                                                .write
		.sgdma_rx_descriptor_write_writedata                   (sgdma_rx_descriptor_write_writedata),                           //                                                .writedata
		.sgdma_rx_m_write_address                              (sgdma_rx_m_write_address),                                      //                                sgdma_rx_m_write.address
		.sgdma_rx_m_write_waitrequest                          (sgdma_rx_m_write_waitrequest),                                  //                                                .waitrequest
		.sgdma_rx_m_write_byteenable                           (sgdma_rx_m_write_byteenable),                                   //                                                .byteenable
		.sgdma_rx_m_write_write                                (sgdma_rx_m_write_write),                                        //                                                .write
		.sgdma_rx_m_write_writedata                            (sgdma_rx_m_write_writedata),                                    //                                                .writedata
		.sgdma_tx_descriptor_read_address                      (sgdma_tx_descriptor_read_address),                              //                        sgdma_tx_descriptor_read.address
		.sgdma_tx_descriptor_read_waitrequest                  (sgdma_tx_descriptor_read_waitrequest),                          //                                                .waitrequest
		.sgdma_tx_descriptor_read_read                         (sgdma_tx_descriptor_read_read),                                 //                                                .read
		.sgdma_tx_descriptor_read_readdata                     (sgdma_tx_descriptor_read_readdata),                             //                                                .readdata
		.sgdma_tx_descriptor_read_readdatavalid                (sgdma_tx_descriptor_read_readdatavalid),                        //                                                .readdatavalid
		.sgdma_tx_descriptor_write_address                     (sgdma_tx_descriptor_write_address),                             //                       sgdma_tx_descriptor_write.address
		.sgdma_tx_descriptor_write_waitrequest                 (sgdma_tx_descriptor_write_waitrequest),                         //                                                .waitrequest
		.sgdma_tx_descriptor_write_write                       (sgdma_tx_descriptor_write_write),                               //                                                .write
		.sgdma_tx_descriptor_write_writedata                   (sgdma_tx_descriptor_write_writedata),                           //                                                .writedata
		.sgdma_tx_m_read_address                               (sgdma_tx_m_read_address),                                       //                                 sgdma_tx_m_read.address
		.sgdma_tx_m_read_waitrequest                           (sgdma_tx_m_read_waitrequest),                                   //                                                .waitrequest
		.sgdma_tx_m_read_read                                  (sgdma_tx_m_read_read),                                          //                                                .read
		.sgdma_tx_m_read_readdata                              (sgdma_tx_m_read_readdata),                                      //                                                .readdata
		.sgdma_tx_m_read_readdatavalid                         (sgdma_tx_m_read_readdatavalid),                                 //                                                .readdatavalid
		.descriptor_memory_s1_address                          (mm_interconnect_0_descriptor_memory_s1_address),                //                            descriptor_memory_s1.address
		.descriptor_memory_s1_write                            (mm_interconnect_0_descriptor_memory_s1_write),                  //                                                .write
		.descriptor_memory_s1_readdata                         (mm_interconnect_0_descriptor_memory_s1_readdata),               //                                                .readdata
		.descriptor_memory_s1_writedata                        (mm_interconnect_0_descriptor_memory_s1_writedata),              //                                                .writedata
		.descriptor_memory_s1_byteenable                       (mm_interconnect_0_descriptor_memory_s1_byteenable),             //                                                .byteenable
		.descriptor_memory_s1_chipselect                       (mm_interconnect_0_descriptor_memory_s1_chipselect),             //                                                .chipselect
		.descriptor_memory_s1_clken                            (mm_interconnect_0_descriptor_memory_s1_clken),                  //                                                .clken
		.mm_clock_crossing_bridge_0_s0_address                 (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_address),       //                   mm_clock_crossing_bridge_0_s0.address
		.mm_clock_crossing_bridge_0_s0_write                   (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_write),         //                                                .write
		.mm_clock_crossing_bridge_0_s0_read                    (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_read),          //                                                .read
		.mm_clock_crossing_bridge_0_s0_readdata                (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdata),      //                                                .readdata
		.mm_clock_crossing_bridge_0_s0_writedata               (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_writedata),     //                                                .writedata
		.mm_clock_crossing_bridge_0_s0_burstcount              (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_burstcount),    //                                                .burstcount
		.mm_clock_crossing_bridge_0_s0_byteenable              (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_byteenable),    //                                                .byteenable
		.mm_clock_crossing_bridge_0_s0_readdatavalid           (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_readdatavalid), //                                                .readdatavalid
		.mm_clock_crossing_bridge_0_s0_waitrequest             (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_waitrequest),   //                                                .waitrequest
		.mm_clock_crossing_bridge_0_s0_debugaccess             (mm_interconnect_0_mm_clock_crossing_bridge_0_s0_debugaccess),   //                                                .debugaccess
		.nios2_gen2_debug_mem_slave_address                    (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),          //                      nios2_gen2_debug_mem_slave.address
		.nios2_gen2_debug_mem_slave_write                      (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),            //                                                .write
		.nios2_gen2_debug_mem_slave_read                       (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),             //                                                .read
		.nios2_gen2_debug_mem_slave_readdata                   (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),         //                                                .readdata
		.nios2_gen2_debug_mem_slave_writedata                  (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),        //                                                .writedata
		.nios2_gen2_debug_mem_slave_byteenable                 (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),       //                                                .byteenable
		.nios2_gen2_debug_mem_slave_waitrequest                (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest),      //                                                .waitrequest
		.nios2_gen2_debug_mem_slave_debugaccess                (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess),      //                                                .debugaccess
		.pll_pll_slave_address                                 (mm_interconnect_0_pll_pll_slave_address),                       //                                   pll_pll_slave.address
		.pll_pll_slave_write                                   (mm_interconnect_0_pll_pll_slave_write),                         //                                                .write
		.pll_pll_slave_read                                    (mm_interconnect_0_pll_pll_slave_read),                          //                                                .read
		.pll_pll_slave_readdata                                (mm_interconnect_0_pll_pll_slave_readdata),                      //                                                .readdata
		.pll_pll_slave_writedata                               (mm_interconnect_0_pll_pll_slave_writedata),                     //                                                .writedata
		.sgdma_rx_csr_address                                  (mm_interconnect_0_sgdma_rx_csr_address),                        //                                    sgdma_rx_csr.address
		.sgdma_rx_csr_write                                    (mm_interconnect_0_sgdma_rx_csr_write),                          //                                                .write
		.sgdma_rx_csr_read                                     (mm_interconnect_0_sgdma_rx_csr_read),                           //                                                .read
		.sgdma_rx_csr_readdata                                 (mm_interconnect_0_sgdma_rx_csr_readdata),                       //                                                .readdata
		.sgdma_rx_csr_writedata                                (mm_interconnect_0_sgdma_rx_csr_writedata),                      //                                                .writedata
		.sgdma_rx_csr_chipselect                               (mm_interconnect_0_sgdma_rx_csr_chipselect),                     //                                                .chipselect
		.sgdma_tx_csr_address                                  (mm_interconnect_0_sgdma_tx_csr_address),                        //                                    sgdma_tx_csr.address
		.sgdma_tx_csr_write                                    (mm_interconnect_0_sgdma_tx_csr_write),                          //                                                .write
		.sgdma_tx_csr_read                                     (mm_interconnect_0_sgdma_tx_csr_read),                           //                                                .read
		.sgdma_tx_csr_readdata                                 (mm_interconnect_0_sgdma_tx_csr_readdata),                       //                                                .readdata
		.sgdma_tx_csr_writedata                                (mm_interconnect_0_sgdma_tx_csr_writedata),                      //                                                .writedata
		.sgdma_tx_csr_chipselect                               (mm_interconnect_0_sgdma_tx_csr_chipselect),                     //                                                .chipselect
		.slow_periph_bridge_s0_address                         (mm_interconnect_0_slow_periph_bridge_s0_address),               //                           slow_periph_bridge_s0.address
		.slow_periph_bridge_s0_write                           (mm_interconnect_0_slow_periph_bridge_s0_write),                 //                                                .write
		.slow_periph_bridge_s0_read                            (mm_interconnect_0_slow_periph_bridge_s0_read),                  //                                                .read
		.slow_periph_bridge_s0_readdata                        (mm_interconnect_0_slow_periph_bridge_s0_readdata),              //                                                .readdata
		.slow_periph_bridge_s0_writedata                       (mm_interconnect_0_slow_periph_bridge_s0_writedata),             //                                                .writedata
		.slow_periph_bridge_s0_burstcount                      (mm_interconnect_0_slow_periph_bridge_s0_burstcount),            //                                                .burstcount
		.slow_periph_bridge_s0_byteenable                      (mm_interconnect_0_slow_periph_bridge_s0_byteenable),            //                                                .byteenable
		.slow_periph_bridge_s0_readdatavalid                   (mm_interconnect_0_slow_periph_bridge_s0_readdatavalid),         //                                                .readdatavalid
		.slow_periph_bridge_s0_waitrequest                     (mm_interconnect_0_slow_periph_bridge_s0_waitrequest),           //                                                .waitrequest
		.slow_periph_bridge_s0_debugaccess                     (mm_interconnect_0_slow_periph_bridge_s0_debugaccess),           //                                                .debugaccess
		.tse_mac_control_port_address                          (mm_interconnect_0_tse_mac_control_port_address),                //                            tse_mac_control_port.address
		.tse_mac_control_port_write                            (mm_interconnect_0_tse_mac_control_port_write),                  //                                                .write
		.tse_mac_control_port_read                             (mm_interconnect_0_tse_mac_control_port_read),                   //                                                .read
		.tse_mac_control_port_readdata                         (mm_interconnect_0_tse_mac_control_port_readdata),               //                                                .readdata
		.tse_mac_control_port_writedata                        (mm_interconnect_0_tse_mac_control_port_writedata),              //                                                .writedata
		.tse_mac_control_port_waitrequest                      (mm_interconnect_0_tse_mac_control_port_waitrequest)             //                                                .waitrequest
	);

	DECA_Qsys_mm_interconnect_1 mm_interconnect_1 (
		.pll_c0_clk                                              (pll_c0_clk),                                                        //                                            pll_c0.clk
		.pll_c2_clk                                              (pll_c2_clk),                                                        //                                            pll_c2.clk
		.jtag_uart_reset_reset_bridge_in_reset_reset             (rst_controller_002_reset_out_reset),                                //             jtag_uart_reset_reset_bridge_in_reset.reset
		.slow_periph_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                                    // slow_periph_bridge_m0_reset_reset_bridge_in_reset.reset
		.slow_periph_bridge_m0_address                           (slow_periph_bridge_m0_address),                                     //                             slow_periph_bridge_m0.address
		.slow_periph_bridge_m0_waitrequest                       (slow_periph_bridge_m0_waitrequest),                                 //                                                  .waitrequest
		.slow_periph_bridge_m0_burstcount                        (slow_periph_bridge_m0_burstcount),                                  //                                                  .burstcount
		.slow_periph_bridge_m0_byteenable                        (slow_periph_bridge_m0_byteenable),                                  //                                                  .byteenable
		.slow_periph_bridge_m0_read                              (slow_periph_bridge_m0_read),                                        //                                                  .read
		.slow_periph_bridge_m0_readdata                          (slow_periph_bridge_m0_readdata),                                    //                                                  .readdata
		.slow_periph_bridge_m0_readdatavalid                     (slow_periph_bridge_m0_readdatavalid),                               //                                                  .readdatavalid
		.slow_periph_bridge_m0_write                             (slow_periph_bridge_m0_write),                                       //                                                  .write
		.slow_periph_bridge_m0_writedata                         (slow_periph_bridge_m0_writedata),                                   //                                                  .writedata
		.slow_periph_bridge_m0_debugaccess                       (slow_periph_bridge_m0_debugaccess),                                 //                                                  .debugaccess
		.ddr3_status_s1_address                                  (mm_interconnect_1_ddr3_status_s1_address),                          //                                    ddr3_status_s1.address
		.ddr3_status_s1_readdata                                 (mm_interconnect_1_ddr3_status_s1_readdata),                         //                                                  .readdata
		.dipsw_pio_s1_address                                    (mm_interconnect_1_dipsw_pio_s1_address),                            //                                      dipsw_pio_s1.address
		.dipsw_pio_s1_write                                      (mm_interconnect_1_dipsw_pio_s1_write),                              //                                                  .write
		.dipsw_pio_s1_readdata                                   (mm_interconnect_1_dipsw_pio_s1_readdata),                           //                                                  .readdata
		.dipsw_pio_s1_writedata                                  (mm_interconnect_1_dipsw_pio_s1_writedata),                          //                                                  .writedata
		.dipsw_pio_s1_chipselect                                 (mm_interconnect_1_dipsw_pio_s1_chipselect),                         //                                                  .chipselect
		.high_res_timer_s1_address                               (mm_interconnect_1_high_res_timer_s1_address),                       //                                 high_res_timer_s1.address
		.high_res_timer_s1_write                                 (mm_interconnect_1_high_res_timer_s1_write),                         //                                                  .write
		.high_res_timer_s1_readdata                              (mm_interconnect_1_high_res_timer_s1_readdata),                      //                                                  .readdata
		.high_res_timer_s1_writedata                             (mm_interconnect_1_high_res_timer_s1_writedata),                     //                                                  .writedata
		.high_res_timer_s1_chipselect                            (mm_interconnect_1_high_res_timer_s1_chipselect),                    //                                                  .chipselect
		.jtag_uart_avalon_jtag_slave_address                     (mm_interconnect_1_jtag_uart_avalon_jtag_slave_address),             //                       jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                       (mm_interconnect_1_jtag_uart_avalon_jtag_slave_write),               //                                                  .write
		.jtag_uart_avalon_jtag_slave_read                        (mm_interconnect_1_jtag_uart_avalon_jtag_slave_read),                //                                                  .read
		.jtag_uart_avalon_jtag_slave_readdata                    (mm_interconnect_1_jtag_uart_avalon_jtag_slave_readdata),            //                                                  .readdata
		.jtag_uart_avalon_jtag_slave_writedata                   (mm_interconnect_1_jtag_uart_avalon_jtag_slave_writedata),           //                                                  .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                 (mm_interconnect_1_jtag_uart_avalon_jtag_slave_waitrequest),         //                                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                  (mm_interconnect_1_jtag_uart_avalon_jtag_slave_chipselect),          //                                                  .chipselect
		.led_pio_s1_address                                      (mm_interconnect_1_led_pio_s1_address),                              //                                        led_pio_s1.address
		.led_pio_s1_write                                        (mm_interconnect_1_led_pio_s1_write),                                //                                                  .write
		.led_pio_s1_readdata                                     (mm_interconnect_1_led_pio_s1_readdata),                             //                                                  .readdata
		.led_pio_s1_writedata                                    (mm_interconnect_1_led_pio_s1_writedata),                            //                                                  .writedata
		.led_pio_s1_chipselect                                   (mm_interconnect_1_led_pio_s1_chipselect),                           //                                                  .chipselect
		.nENET_reg_reset_s1_address                              (mm_interconnect_1_nenet_reg_reset_s1_address),                      //                                nENET_reg_reset_s1.address
		.nENET_reg_reset_s1_write                                (mm_interconnect_1_nenet_reg_reset_s1_write),                        //                                                  .write
		.nENET_reg_reset_s1_readdata                             (mm_interconnect_1_nenet_reg_reset_s1_readdata),                     //                                                  .readdata
		.nENET_reg_reset_s1_writedata                            (mm_interconnect_1_nenet_reg_reset_s1_writedata),                    //                                                  .writedata
		.nENET_reg_reset_s1_chipselect                           (mm_interconnect_1_nenet_reg_reset_s1_chipselect),                   //                                                  .chipselect
		.performance_counter_control_slave_address               (mm_interconnect_1_performance_counter_control_slave_address),       //                 performance_counter_control_slave.address
		.performance_counter_control_slave_write                 (mm_interconnect_1_performance_counter_control_slave_write),         //                                                  .write
		.performance_counter_control_slave_readdata              (mm_interconnect_1_performance_counter_control_slave_readdata),      //                                                  .readdata
		.performance_counter_control_slave_writedata             (mm_interconnect_1_performance_counter_control_slave_writedata),     //                                                  .writedata
		.performance_counter_control_slave_begintransfer         (mm_interconnect_1_performance_counter_control_slave_begintransfer), //                                                  .begintransfer
		.sys_timer_s1_address                                    (mm_interconnect_1_sys_timer_s1_address),                            //                                      sys_timer_s1.address
		.sys_timer_s1_write                                      (mm_interconnect_1_sys_timer_s1_write),                              //                                                  .write
		.sys_timer_s1_readdata                                   (mm_interconnect_1_sys_timer_s1_readdata),                           //                                                  .readdata
		.sys_timer_s1_writedata                                  (mm_interconnect_1_sys_timer_s1_writedata),                          //                                                  .writedata
		.sys_timer_s1_chipselect                                 (mm_interconnect_1_sys_timer_s1_chipselect),                         //                                                  .chipselect
		.sysid_control_slave_address                             (mm_interconnect_1_sysid_control_slave_address),                     //                               sysid_control_slave.address
		.sysid_control_slave_readdata                            (mm_interconnect_1_sysid_control_slave_readdata),                    //                                                  .readdata
		.user_pio_pushbtn_s1_address                             (mm_interconnect_1_user_pio_pushbtn_s1_address),                     //                               user_pio_pushbtn_s1.address
		.user_pio_pushbtn_s1_readdata                            (mm_interconnect_1_user_pio_pushbtn_s1_readdata)                     //                                                  .readdata
	);

	DECA_Qsys_mm_interconnect_2 mm_interconnect_2 (
		.mem_if_ddr3_emif_afi_clk_clk                                    (mem_if_ddr3_emif_afi_clk_clk),                              //                                  mem_if_ddr3_emif_afi_clk.clk
		.mem_if_ddr3_emif_soft_reset_reset_bridge_in_reset_reset         (rst_controller_005_reset_out_reset),                        //         mem_if_ddr3_emif_soft_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset (rst_controller_005_reset_out_reset),                        // mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_0_m0_address                           (mm_clock_crossing_bridge_0_m0_address),                     //                             mm_clock_crossing_bridge_0_m0.address
		.mm_clock_crossing_bridge_0_m0_waitrequest                       (mm_clock_crossing_bridge_0_m0_waitrequest),                 //                                                          .waitrequest
		.mm_clock_crossing_bridge_0_m0_burstcount                        (mm_clock_crossing_bridge_0_m0_burstcount),                  //                                                          .burstcount
		.mm_clock_crossing_bridge_0_m0_byteenable                        (mm_clock_crossing_bridge_0_m0_byteenable),                  //                                                          .byteenable
		.mm_clock_crossing_bridge_0_m0_read                              (mm_clock_crossing_bridge_0_m0_read),                        //                                                          .read
		.mm_clock_crossing_bridge_0_m0_readdata                          (mm_clock_crossing_bridge_0_m0_readdata),                    //                                                          .readdata
		.mm_clock_crossing_bridge_0_m0_readdatavalid                     (mm_clock_crossing_bridge_0_m0_readdatavalid),               //                                                          .readdatavalid
		.mm_clock_crossing_bridge_0_m0_write                             (mm_clock_crossing_bridge_0_m0_write),                       //                                                          .write
		.mm_clock_crossing_bridge_0_m0_writedata                         (mm_clock_crossing_bridge_0_m0_writedata),                   //                                                          .writedata
		.mm_clock_crossing_bridge_0_m0_debugaccess                       (mm_clock_crossing_bridge_0_m0_debugaccess),                 //                                                          .debugaccess
		.mem_if_ddr3_emif_avl_address                                    (mm_interconnect_2_mem_if_ddr3_emif_avl_address),            //                                      mem_if_ddr3_emif_avl.address
		.mem_if_ddr3_emif_avl_write                                      (mm_interconnect_2_mem_if_ddr3_emif_avl_write),              //                                                          .write
		.mem_if_ddr3_emif_avl_read                                       (mm_interconnect_2_mem_if_ddr3_emif_avl_read),               //                                                          .read
		.mem_if_ddr3_emif_avl_readdata                                   (mm_interconnect_2_mem_if_ddr3_emif_avl_readdata),           //                                                          .readdata
		.mem_if_ddr3_emif_avl_writedata                                  (mm_interconnect_2_mem_if_ddr3_emif_avl_writedata),          //                                                          .writedata
		.mem_if_ddr3_emif_avl_beginbursttransfer                         (mm_interconnect_2_mem_if_ddr3_emif_avl_beginbursttransfer), //                                                          .beginbursttransfer
		.mem_if_ddr3_emif_avl_burstcount                                 (mm_interconnect_2_mem_if_ddr3_emif_avl_burstcount),         //                                                          .burstcount
		.mem_if_ddr3_emif_avl_byteenable                                 (mm_interconnect_2_mem_if_ddr3_emif_avl_byteenable),         //                                                          .byteenable
		.mem_if_ddr3_emif_avl_readdatavalid                              (mm_interconnect_2_mem_if_ddr3_emif_avl_readdatavalid),      //                                                          .readdatavalid
		.mem_if_ddr3_emif_avl_waitrequest                                (~mm_interconnect_2_mem_if_ddr3_emif_avl_waitrequest)        //                                                          .waitrequest
	);

	DECA_Qsys_irq_mapper irq_mapper (
		.clk           (pll_c0_clk),                         //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (nios2_gen2_irq_irq)                  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_c2_clk),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (pll_c2_clk),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_clk),                         //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	DECA_Qsys_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (6),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (pll_c0_clk),                            // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_001_reset_out_reset),    // in_rst_0.reset
		.in_0_data           (tse_mac_receive_data),                  //     in_0.data
		.in_0_valid          (tse_mac_receive_valid),                 //         .valid
		.in_0_ready          (tse_mac_receive_ready),                 //         .ready
		.in_0_startofpacket  (tse_mac_receive_startofpacket),         //         .startofpacket
		.in_0_endofpacket    (tse_mac_receive_endofpacket),           //         .endofpacket
		.in_0_empty          (tse_mac_receive_empty),                 //         .empty
		.in_0_error          (tse_mac_receive_error),                 //         .error
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_out_0_error)          //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (pll_c2_clk),                     //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (pll_c0_clk),                             //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset),   // reset_in1.reset
		.clk            (pll_c0_clk),                             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset), // reset_in1.reset
		.clk            (),                                     //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset), // reset_in1.reset
		.clk            (),                                     //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset), // reset_in1.reset
		.clk            (mem_if_ddr3_emif_afi_clk_clk),         //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
