// usb20sr_refdes.v

// Generated using ACDS version 15.0 139

`timescale 1 ps / 1 ps
module usb20sr_refdes (
		input  wire       altpll_0_areset_conduit_export,      //      altpll_0_areset_conduit.export
		output wire       altpll_0_locked_conduit_export,      //      altpll_0_locked_conduit.export
		output wire       altpll_0_phasedone_conduit_export,   //   altpll_0_phasedone_conduit.export
		input  wire       osc_clk_clk,                         //                      osc_clk.clk
		input  wire       reset_reset_n,                       //                        reset.reset_n
		output wire       rst_pio_external_connection_export,  //  rst_pio_external_connection.export
		input  wire       u20_clk_out_clk,                     //                  u20_clk_out.clk
		inout  wire [7:0] usb20sr_conduit_end_Data,            //          usb20sr_conduit_end.Data
		output wire       usb20sr_conduit_end_Stp,             //                             .Stp
		input  wire       usb20sr_conduit_end_Dir,             //                             .Dir
		input  wire       usb20sr_conduit_end_Nxt,             //                             .Nxt
		input  wire       usb20sr_conduit_end_phy_clk,         //                             .phy_clk
		output wire       usb20sr_conduit_end_phy_reset_n,     //                             .phy_reset_n
		output wire       usb20sr_conduit_end_phy_cs_n,        //                             .phy_cs_n
		input  wire       usb20sr_conduit_end_Ext_reset_in,    //                             .Ext_reset_in
		output wire [7:0] user_led_external_connection_export  // user_led_external_connection.export
	);

	wire         altpll_0_c0_clk;                                              // altpll_0:c0 -> [ccb_slow_per:s0_clk, ccb_usb:s0_clk, dma_0:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, jtag_uart_0:clk, mm_interconnect_0:altpll_0_c0_clk, nios2_qsys_0:clk, onchip_memory:clk, rst_controller_002:clk, rst_controller_004:clk]
	wire         altpll_0_c2_clk;                                              // altpll_0:c2 -> [ccb_slow_per:m0_clk, irq_synchronizer:receiver_clk, mm_interconnect_2:altpll_0_c2_clk, rst_controller_001:clk, rst_pio:clk, timer_0:clk, user_led:clk]
	wire  [31:0] nios2_qsys_0_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                         // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [25:0] nios2_qsys_0_data_master_address;                             // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                          // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_readdatavalid;                       // mm_interconnect_0:nios2_qsys_0_data_master_readdatavalid -> nios2_qsys_0:d_readdatavalid
	wire         nios2_qsys_0_data_master_write;                               // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                           // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [24:0] nios2_qsys_0_instruction_master_address;                      // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                         // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         nios2_qsys_0_instruction_master_readdatavalid;                // mm_interconnect_0:nios2_qsys_0_instruction_master_readdatavalid -> nios2_qsys_0:i_readdatavalid
	wire         dma_0_read_master_chipselect;                                 // dma_0:read_chipselect -> mm_interconnect_0:dma_0_read_master_chipselect
	wire  [31:0] dma_0_read_master_readdata;                                   // mm_interconnect_0:dma_0_read_master_readdata -> dma_0:read_readdata
	wire         dma_0_read_master_waitrequest;                                // mm_interconnect_0:dma_0_read_master_waitrequest -> dma_0:read_waitrequest
	wire  [24:0] dma_0_read_master_address;                                    // dma_0:read_address -> mm_interconnect_0:dma_0_read_master_address
	wire         dma_0_read_master_read;                                       // dma_0:read_read_n -> mm_interconnect_0:dma_0_read_master_read
	wire         dma_0_read_master_readdatavalid;                              // mm_interconnect_0:dma_0_read_master_readdatavalid -> dma_0:read_readdatavalid
	wire         dma_0_write_master_chipselect;                                // dma_0:write_chipselect -> mm_interconnect_0:dma_0_write_master_chipselect
	wire         dma_0_write_master_waitrequest;                               // mm_interconnect_0:dma_0_write_master_waitrequest -> dma_0:write_waitrequest
	wire  [24:0] dma_0_write_master_address;                                   // dma_0:write_address -> mm_interconnect_0:dma_0_write_master_address
	wire   [3:0] dma_0_write_master_byteenable;                                // dma_0:write_byteenable -> mm_interconnect_0:dma_0_write_master_byteenable
	wire         dma_0_write_master_write;                                     // dma_0:write_write_n -> mm_interconnect_0:dma_0_write_master_write
	wire  [31:0] dma_0_write_master_writedata;                                 // dma_0:write_writedata -> mm_interconnect_0:dma_0_write_master_writedata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire         mm_interconnect_0_dma_0_control_port_slave_chipselect;        // mm_interconnect_0:dma_0_control_port_slave_chipselect -> dma_0:dma_ctl_chipselect
	wire  [24:0] mm_interconnect_0_dma_0_control_port_slave_readdata;          // dma_0:dma_ctl_readdata -> mm_interconnect_0:dma_0_control_port_slave_readdata
	wire   [2:0] mm_interconnect_0_dma_0_control_port_slave_address;           // mm_interconnect_0:dma_0_control_port_slave_address -> dma_0:dma_ctl_address
	wire         mm_interconnect_0_dma_0_control_port_slave_write;             // mm_interconnect_0:dma_0_control_port_slave_write -> dma_0:dma_ctl_write_n
	wire  [24:0] mm_interconnect_0_dma_0_control_port_slave_writedata;         // mm_interconnect_0:dma_0_control_port_slave_writedata -> dma_0:dma_ctl_writedata
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;    // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest; // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;                // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                 // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                    // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                   // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;               // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire  [31:0] mm_interconnect_0_ccb_usb_s0_readdata;                        // ccb_usb:s0_readdata -> mm_interconnect_0:ccb_usb_s0_readdata
	wire         mm_interconnect_0_ccb_usb_s0_waitrequest;                     // ccb_usb:s0_waitrequest -> mm_interconnect_0:ccb_usb_s0_waitrequest
	wire         mm_interconnect_0_ccb_usb_s0_debugaccess;                     // mm_interconnect_0:ccb_usb_s0_debugaccess -> ccb_usb:s0_debugaccess
	wire  [20:0] mm_interconnect_0_ccb_usb_s0_address;                         // mm_interconnect_0:ccb_usb_s0_address -> ccb_usb:s0_address
	wire         mm_interconnect_0_ccb_usb_s0_read;                            // mm_interconnect_0:ccb_usb_s0_read -> ccb_usb:s0_read
	wire   [3:0] mm_interconnect_0_ccb_usb_s0_byteenable;                      // mm_interconnect_0:ccb_usb_s0_byteenable -> ccb_usb:s0_byteenable
	wire         mm_interconnect_0_ccb_usb_s0_readdatavalid;                   // ccb_usb:s0_readdatavalid -> mm_interconnect_0:ccb_usb_s0_readdatavalid
	wire         mm_interconnect_0_ccb_usb_s0_write;                           // mm_interconnect_0:ccb_usb_s0_write -> ccb_usb:s0_write
	wire  [31:0] mm_interconnect_0_ccb_usb_s0_writedata;                       // mm_interconnect_0:ccb_usb_s0_writedata -> ccb_usb:s0_writedata
	wire   [0:0] mm_interconnect_0_ccb_usb_s0_burstcount;                      // mm_interconnect_0:ccb_usb_s0_burstcount -> ccb_usb:s0_burstcount
	wire  [31:0] mm_interconnect_0_ccb_slow_per_s0_readdata;                   // ccb_slow_per:s0_readdata -> mm_interconnect_0:ccb_slow_per_s0_readdata
	wire         mm_interconnect_0_ccb_slow_per_s0_waitrequest;                // ccb_slow_per:s0_waitrequest -> mm_interconnect_0:ccb_slow_per_s0_waitrequest
	wire         mm_interconnect_0_ccb_slow_per_s0_debugaccess;                // mm_interconnect_0:ccb_slow_per_s0_debugaccess -> ccb_slow_per:s0_debugaccess
	wire   [6:0] mm_interconnect_0_ccb_slow_per_s0_address;                    // mm_interconnect_0:ccb_slow_per_s0_address -> ccb_slow_per:s0_address
	wire         mm_interconnect_0_ccb_slow_per_s0_read;                       // mm_interconnect_0:ccb_slow_per_s0_read -> ccb_slow_per:s0_read
	wire   [3:0] mm_interconnect_0_ccb_slow_per_s0_byteenable;                 // mm_interconnect_0:ccb_slow_per_s0_byteenable -> ccb_slow_per:s0_byteenable
	wire         mm_interconnect_0_ccb_slow_per_s0_readdatavalid;              // ccb_slow_per:s0_readdatavalid -> mm_interconnect_0:ccb_slow_per_s0_readdatavalid
	wire         mm_interconnect_0_ccb_slow_per_s0_write;                      // mm_interconnect_0:ccb_slow_per_s0_write -> ccb_slow_per:s0_write
	wire  [31:0] mm_interconnect_0_ccb_slow_per_s0_writedata;                  // mm_interconnect_0:ccb_slow_per_s0_writedata -> ccb_slow_per:s0_writedata
	wire   [0:0] mm_interconnect_0_ccb_slow_per_s0_burstcount;                 // mm_interconnect_0:ccb_slow_per_s0_burstcount -> ccb_slow_per:s0_burstcount
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                  // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory_s1_address;                   // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                     // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                 // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                     // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_onchip_memory_s2_chipselect;                // mm_interconnect_0:onchip_memory_s2_chipselect -> onchip_memory:chipselect2
	wire  [31:0] mm_interconnect_0_onchip_memory_s2_readdata;                  // onchip_memory:readdata2 -> mm_interconnect_0:onchip_memory_s2_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory_s2_address;                   // mm_interconnect_0:onchip_memory_s2_address -> onchip_memory:address2
	wire   [3:0] mm_interconnect_0_onchip_memory_s2_byteenable;                // mm_interconnect_0:onchip_memory_s2_byteenable -> onchip_memory:byteenable2
	wire         mm_interconnect_0_onchip_memory_s2_write;                     // mm_interconnect_0:onchip_memory_s2_write -> onchip_memory:write2
	wire  [31:0] mm_interconnect_0_onchip_memory_s2_writedata;                 // mm_interconnect_0:onchip_memory_s2_writedata -> onchip_memory:writedata2
	wire         mm_interconnect_0_onchip_memory_s2_clken;                     // mm_interconnect_0:onchip_memory_s2_clken -> onchip_memory:clken2
	wire         ccb_usb_m0_waitrequest;                                       // mm_interconnect_1:ccb_usb_m0_waitrequest -> ccb_usb:m0_waitrequest
	wire  [31:0] ccb_usb_m0_readdata;                                          // mm_interconnect_1:ccb_usb_m0_readdata -> ccb_usb:m0_readdata
	wire         ccb_usb_m0_debugaccess;                                       // ccb_usb:m0_debugaccess -> mm_interconnect_1:ccb_usb_m0_debugaccess
	wire  [20:0] ccb_usb_m0_address;                                           // ccb_usb:m0_address -> mm_interconnect_1:ccb_usb_m0_address
	wire         ccb_usb_m0_read;                                              // ccb_usb:m0_read -> mm_interconnect_1:ccb_usb_m0_read
	wire   [3:0] ccb_usb_m0_byteenable;                                        // ccb_usb:m0_byteenable -> mm_interconnect_1:ccb_usb_m0_byteenable
	wire         ccb_usb_m0_readdatavalid;                                     // mm_interconnect_1:ccb_usb_m0_readdatavalid -> ccb_usb:m0_readdatavalid
	wire  [31:0] ccb_usb_m0_writedata;                                         // ccb_usb:m0_writedata -> mm_interconnect_1:ccb_usb_m0_writedata
	wire         ccb_usb_m0_write;                                             // ccb_usb:m0_write -> mm_interconnect_1:ccb_usb_m0_write
	wire   [0:0] ccb_usb_m0_burstcount;                                        // ccb_usb:m0_burstcount -> mm_interconnect_1:ccb_usb_m0_burstcount
	wire         mm_interconnect_1_usb20sr_avalon_slave_0_chipselect;          // mm_interconnect_1:usb20sr_avalon_slave_0_chipselect -> usb20sr:chipselect
	wire  [31:0] mm_interconnect_1_usb20sr_avalon_slave_0_readdata;            // usb20sr:readdata -> mm_interconnect_1:usb20sr_avalon_slave_0_readdata
	wire         mm_interconnect_1_usb20sr_avalon_slave_0_waitrequest;         // usb20sr:waitrequest -> mm_interconnect_1:usb20sr_avalon_slave_0_waitrequest
	wire  [18:0] mm_interconnect_1_usb20sr_avalon_slave_0_address;             // mm_interconnect_1:usb20sr_avalon_slave_0_address -> usb20sr:address
	wire         mm_interconnect_1_usb20sr_avalon_slave_0_read;                // mm_interconnect_1:usb20sr_avalon_slave_0_read -> usb20sr:read_n
	wire   [3:0] mm_interconnect_1_usb20sr_avalon_slave_0_byteenable;          // mm_interconnect_1:usb20sr_avalon_slave_0_byteenable -> usb20sr:byteenable_n
	wire         mm_interconnect_1_usb20sr_avalon_slave_0_readdatavalid;       // usb20sr:readdatavalid -> mm_interconnect_1:usb20sr_avalon_slave_0_readdatavalid
	wire         mm_interconnect_1_usb20sr_avalon_slave_0_write;               // mm_interconnect_1:usb20sr_avalon_slave_0_write -> usb20sr:write_n
	wire  [31:0] mm_interconnect_1_usb20sr_avalon_slave_0_writedata;           // mm_interconnect_1:usb20sr_avalon_slave_0_writedata -> usb20sr:writedata
	wire         ccb_slow_per_m0_waitrequest;                                  // mm_interconnect_2:ccb_slow_per_m0_waitrequest -> ccb_slow_per:m0_waitrequest
	wire  [31:0] ccb_slow_per_m0_readdata;                                     // mm_interconnect_2:ccb_slow_per_m0_readdata -> ccb_slow_per:m0_readdata
	wire         ccb_slow_per_m0_debugaccess;                                  // ccb_slow_per:m0_debugaccess -> mm_interconnect_2:ccb_slow_per_m0_debugaccess
	wire   [6:0] ccb_slow_per_m0_address;                                      // ccb_slow_per:m0_address -> mm_interconnect_2:ccb_slow_per_m0_address
	wire         ccb_slow_per_m0_read;                                         // ccb_slow_per:m0_read -> mm_interconnect_2:ccb_slow_per_m0_read
	wire   [3:0] ccb_slow_per_m0_byteenable;                                   // ccb_slow_per:m0_byteenable -> mm_interconnect_2:ccb_slow_per_m0_byteenable
	wire         ccb_slow_per_m0_readdatavalid;                                // mm_interconnect_2:ccb_slow_per_m0_readdatavalid -> ccb_slow_per:m0_readdatavalid
	wire  [31:0] ccb_slow_per_m0_writedata;                                    // ccb_slow_per:m0_writedata -> mm_interconnect_2:ccb_slow_per_m0_writedata
	wire         ccb_slow_per_m0_write;                                        // ccb_slow_per:m0_write -> mm_interconnect_2:ccb_slow_per_m0_write
	wire   [0:0] ccb_slow_per_m0_burstcount;                                   // ccb_slow_per:m0_burstcount -> mm_interconnect_2:ccb_slow_per_m0_burstcount
	wire         mm_interconnect_2_timer_0_s1_chipselect;                      // mm_interconnect_2:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_2_timer_0_s1_readdata;                        // timer_0:readdata -> mm_interconnect_2:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_2_timer_0_s1_address;                         // mm_interconnect_2:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_2_timer_0_s1_write;                           // mm_interconnect_2:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_2_timer_0_s1_writedata;                       // mm_interconnect_2:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_2_user_led_s1_chipselect;                     // mm_interconnect_2:user_led_s1_chipselect -> user_led:chipselect
	wire  [31:0] mm_interconnect_2_user_led_s1_readdata;                       // user_led:readdata -> mm_interconnect_2:user_led_s1_readdata
	wire   [1:0] mm_interconnect_2_user_led_s1_address;                        // mm_interconnect_2:user_led_s1_address -> user_led:address
	wire         mm_interconnect_2_user_led_s1_write;                          // mm_interconnect_2:user_led_s1_write -> user_led:write_n
	wire  [31:0] mm_interconnect_2_user_led_s1_writedata;                      // mm_interconnect_2:user_led_s1_writedata -> user_led:writedata
	wire         mm_interconnect_2_rst_pio_s1_chipselect;                      // mm_interconnect_2:rst_pio_s1_chipselect -> rst_pio:chipselect
	wire  [31:0] mm_interconnect_2_rst_pio_s1_readdata;                        // rst_pio:readdata -> mm_interconnect_2:rst_pio_s1_readdata
	wire   [1:0] mm_interconnect_2_rst_pio_s1_address;                         // mm_interconnect_2:rst_pio_s1_address -> rst_pio:address
	wire         mm_interconnect_2_rst_pio_s1_write;                           // mm_interconnect_2:rst_pio_s1_write -> rst_pio:write_n
	wire  [31:0] mm_interconnect_2_rst_pio_s1_writedata;                       // mm_interconnect_2:rst_pio_s1_writedata -> rst_pio:writedata
	wire         irq_mapper_receiver0_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver2_irq;                                     // dma_0:dma_ctl_irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         irq_mapper_receiver1_irq;                                     // irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                // timer_0:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver3_irq;                                     // irq_synchronizer_001:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                            // usb20sr:irq -> irq_synchronizer_001:receiver_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                           // rst_controller_001:reset_out -> [ccb_slow_per:m0_reset, irq_synchronizer:receiver_reset, mm_interconnect_2:ccb_slow_per_m0_reset_reset_bridge_in_reset_reset, rst_pio:reset_n, timer_0:reset_n, user_led:reset_n]
	wire         rst_controller_002_reset_out_reset;                           // rst_controller_002:reset_out -> [ccb_slow_per:s0_reset, ccb_usb:s0_reset, dma_0:system_reset_n, jtag_uart_0:rst_n, mm_interconnect_0:dma_0_reset_reset_bridge_in_reset_reset, onchip_memory:reset, rst_translator:in_reset]
	wire         rst_controller_002_reset_out_reset_req;                       // rst_controller_002:reset_req -> [onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_003_reset_out_reset;                           // rst_controller_003:reset_out -> [ccb_usb:m0_reset, mm_interconnect_1:ccb_usb_m0_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_004_reset_out_reset;                           // rst_controller_004:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, rst_translator_001:in_reset]
	wire         rst_controller_004_reset_out_reset_req;                       // rst_controller_004:reset_req -> [nios2_qsys_0:reset_req, rst_translator_001:reset_req_in]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                   // nios2_qsys_0:jtag_debug_module_resetrequest -> rst_controller_004:reset_in1
	wire         rst_controller_005_reset_out_reset;                           // rst_controller_005:reset_out -> [irq_synchronizer_001:receiver_reset, mm_interconnect_1:usb20sr_clock_reset_reset_bridge_in_reset_reset, usb20sr:reset_n]

	usb20sr_refdes_altpll_0 altpll_0 (
		.clk       (osc_clk_clk),                                    //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),                 // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0        (altpll_0_c0_clk),                                //                    c0.clk
		.c1        (),                                               //                    c1.clk
		.c2        (altpll_0_c2_clk),                                //                    c2.clk
		.areset    (altpll_0_areset_conduit_export),                 //        areset_conduit.export
		.locked    (altpll_0_locked_conduit_export),                 //        locked_conduit.export
		.phasedone (altpll_0_phasedone_conduit_export)               //     phasedone_conduit.export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (7),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (32),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) ccb_slow_per (
		.m0_clk           (altpll_0_c2_clk),                                 //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),              // m0_reset.reset
		.s0_clk           (altpll_0_c0_clk),                                 //   s0_clk.clk
		.s0_reset         (rst_controller_002_reset_out_reset),              // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_ccb_slow_per_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_ccb_slow_per_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_ccb_slow_per_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_ccb_slow_per_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_ccb_slow_per_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_ccb_slow_per_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_ccb_slow_per_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_ccb_slow_per_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_ccb_slow_per_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_ccb_slow_per_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (ccb_slow_per_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (ccb_slow_per_m0_readdata),                        //         .readdata
		.m0_readdatavalid (ccb_slow_per_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (ccb_slow_per_m0_burstcount),                      //         .burstcount
		.m0_writedata     (ccb_slow_per_m0_writedata),                       //         .writedata
		.m0_address       (ccb_slow_per_m0_address),                         //         .address
		.m0_write         (ccb_slow_per_m0_write),                           //         .write
		.m0_read          (ccb_slow_per_m0_read),                            //         .read
		.m0_byteenable    (ccb_slow_per_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (ccb_slow_per_m0_debugaccess)                      //         .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (21),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (16),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) ccb_usb (
		.m0_clk           (u20_clk_out_clk),                            //   m0_clk.clk
		.m0_reset         (rst_controller_003_reset_out_reset),         // m0_reset.reset
		.s0_clk           (altpll_0_c0_clk),                            //   s0_clk.clk
		.s0_reset         (rst_controller_002_reset_out_reset),         // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_ccb_usb_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_ccb_usb_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_ccb_usb_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_ccb_usb_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_ccb_usb_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_ccb_usb_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_ccb_usb_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_ccb_usb_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_ccb_usb_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_ccb_usb_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (ccb_usb_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (ccb_usb_m0_readdata),                        //         .readdata
		.m0_readdatavalid (ccb_usb_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (ccb_usb_m0_burstcount),                      //         .burstcount
		.m0_writedata     (ccb_usb_m0_writedata),                       //         .writedata
		.m0_address       (ccb_usb_m0_address),                         //         .address
		.m0_write         (ccb_usb_m0_write),                           //         .write
		.m0_read          (ccb_usb_m0_read),                            //         .read
		.m0_byteenable    (ccb_usb_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (ccb_usb_m0_debugaccess)                      //         .debugaccess
	);

	usb20sr_refdes_dma_0 dma_0 (
		.clk                (altpll_0_c0_clk),                                       //                clk.clk
		.system_reset_n     (~rst_controller_002_reset_out_reset),                   //              reset.reset_n
		.dma_ctl_address    (mm_interconnect_0_dma_0_control_port_slave_address),    // control_port_slave.address
		.dma_ctl_chipselect (mm_interconnect_0_dma_0_control_port_slave_chipselect), //                   .chipselect
		.dma_ctl_readdata   (mm_interconnect_0_dma_0_control_port_slave_readdata),   //                   .readdata
		.dma_ctl_write_n    (~mm_interconnect_0_dma_0_control_port_slave_write),     //                   .write_n
		.dma_ctl_writedata  (mm_interconnect_0_dma_0_control_port_slave_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_mapper_receiver2_irq),                              //                irq.irq
		.read_address       (dma_0_read_master_address),                             //        read_master.address
		.read_chipselect    (dma_0_read_master_chipselect),                          //                   .chipselect
		.read_read_n        (dma_0_read_master_read),                                //                   .read_n
		.read_readdata      (dma_0_read_master_readdata),                            //                   .readdata
		.read_readdatavalid (dma_0_read_master_readdatavalid),                       //                   .readdatavalid
		.read_waitrequest   (dma_0_read_master_waitrequest),                         //                   .waitrequest
		.write_address      (dma_0_write_master_address),                            //       write_master.address
		.write_chipselect   (dma_0_write_master_chipselect),                         //                   .chipselect
		.write_waitrequest  (dma_0_write_master_waitrequest),                        //                   .waitrequest
		.write_write_n      (dma_0_write_master_write),                              //                   .write_n
		.write_writedata    (dma_0_write_master_writedata),                          //                   .writedata
		.write_byteenable   (dma_0_write_master_byteenable)                          //                   .byteenable
	);

	usb20sr_refdes_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_0_c0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	usb20sr_refdes_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (altpll_0_c0_clk),                                              //                       clk.clk
		.reset_n                               (~rst_controller_004_reset_out_reset),                          //                   reset_n.reset_n
		.reset_req                             (rst_controller_004_reset_out_reset_req),                       //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_qsys_0_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_0_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	usb20sr_refdes_onchip_memory onchip_memory (
		.address     (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.address2    (mm_interconnect_0_onchip_memory_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_memory_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_memory_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_memory_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_memory_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_memory_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_onchip_memory_s2_byteenable), //       .byteenable
		.clk         (altpll_0_c0_clk),                               //   clk1.clk
		.reset       (rst_controller_002_reset_out_reset),            // reset1.reset
		.reset_req   (rst_controller_002_reset_out_reset_req)         //       .reset_req
	);

	usb20sr_refdes_rst_pio rst_pio (
		.clk        (altpll_0_c2_clk),                         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_2_rst_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_rst_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_rst_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_rst_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_rst_pio_s1_readdata),   //                    .readdata
		.out_port   (rst_pio_external_connection_export)       // external_connection.export
	);

	usb20sr_refdes_timer_0 timer_0 (
		.clk        (altpll_0_c2_clk),                         //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_2_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_2_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_2_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_2_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_2_timer_0_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)            //   irq.irq
	);

	sls_avalon_usb20sr #(
		.IN_DEPTH       (512),
		.OUT_DEPTH      (512),
		.IN_ADR_WIDTH   (9),
		.OUT_ADR_WIDTH  (9),
		.Simulation     (1),
		.Interface_sel  (0),
		.Enum_data_file ("Enum_ram.hex")
	) usb20sr (
		.clk           (u20_clk_out_clk),                                        //          clock.clk
		.reset_n       (~rst_controller_005_reset_out_reset),                    //    clock_reset.reset_n
		.address       (mm_interconnect_1_usb20sr_avalon_slave_0_address),       // avalon_slave_0.address
		.writedata     (mm_interconnect_1_usb20sr_avalon_slave_0_writedata),     //               .writedata
		.chipselect    (mm_interconnect_1_usb20sr_avalon_slave_0_chipselect),    //               .chipselect
		.write_n       (~mm_interconnect_1_usb20sr_avalon_slave_0_write),        //               .write_n
		.read_n        (~mm_interconnect_1_usb20sr_avalon_slave_0_read),         //               .read_n
		.byteenable_n  (~mm_interconnect_1_usb20sr_avalon_slave_0_byteenable),   //               .byteenable_n
		.readdata      (mm_interconnect_1_usb20sr_avalon_slave_0_readdata),      //               .readdata
		.waitrequest   (mm_interconnect_1_usb20sr_avalon_slave_0_waitrequest),   //               .waitrequest
		.readdatavalid (mm_interconnect_1_usb20sr_avalon_slave_0_readdatavalid), //               .readdatavalid
		.irq           (irq_synchronizer_001_receiver_irq),                      //           irq0.irq
		.Data          (usb20sr_conduit_end_Data),                               //    conduit_end.export
		.Stp           (usb20sr_conduit_end_Stp),                                //               .export
		.Dir           (usb20sr_conduit_end_Dir),                                //               .export
		.Nxt           (usb20sr_conduit_end_Nxt),                                //               .export
		.phy_clk       (usb20sr_conduit_end_phy_clk),                            //               .export
		.phy_reset_n   (usb20sr_conduit_end_phy_reset_n),                        //               .export
		.phy_cs_n      (usb20sr_conduit_end_phy_cs_n),                           //               .export
		.Ext_reset_in  (usb20sr_conduit_end_Ext_reset_in)                        //               .export
	);

	usb20sr_refdes_user_led user_led (
		.clk        (altpll_0_c2_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_2_user_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_2_user_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_2_user_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_2_user_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_2_user_led_s1_readdata),   //                    .readdata
		.out_port   (user_led_external_connection_export)       // external_connection.export
	);

	usb20sr_refdes_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                                            (altpll_0_c0_clk),                                              //                                          altpll_0_c0.clk
		.osc_clk_clk_clk                                            (osc_clk_clk),                                                  //                                          osc_clk_clk.clk
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                               // altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.dma_0_reset_reset_bridge_in_reset_reset                    (rst_controller_002_reset_out_reset),                           //                    dma_0_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset           (rst_controller_004_reset_out_reset),                           //           nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.dma_0_read_master_address                                  (dma_0_read_master_address),                                    //                                    dma_0_read_master.address
		.dma_0_read_master_waitrequest                              (dma_0_read_master_waitrequest),                                //                                                     .waitrequest
		.dma_0_read_master_chipselect                               (dma_0_read_master_chipselect),                                 //                                                     .chipselect
		.dma_0_read_master_read                                     (~dma_0_read_master_read),                                      //                                                     .read
		.dma_0_read_master_readdata                                 (dma_0_read_master_readdata),                                   //                                                     .readdata
		.dma_0_read_master_readdatavalid                            (dma_0_read_master_readdatavalid),                              //                                                     .readdatavalid
		.dma_0_write_master_address                                 (dma_0_write_master_address),                                   //                                   dma_0_write_master.address
		.dma_0_write_master_waitrequest                             (dma_0_write_master_waitrequest),                               //                                                     .waitrequest
		.dma_0_write_master_byteenable                              (dma_0_write_master_byteenable),                                //                                                     .byteenable
		.dma_0_write_master_chipselect                              (dma_0_write_master_chipselect),                                //                                                     .chipselect
		.dma_0_write_master_write                                   (~dma_0_write_master_write),                                    //                                                     .write
		.dma_0_write_master_writedata                               (dma_0_write_master_writedata),                                 //                                                     .writedata
		.nios2_qsys_0_data_master_address                           (nios2_qsys_0_data_master_address),                             //                             nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest                       (nios2_qsys_0_data_master_waitrequest),                         //                                                     .waitrequest
		.nios2_qsys_0_data_master_byteenable                        (nios2_qsys_0_data_master_byteenable),                          //                                                     .byteenable
		.nios2_qsys_0_data_master_read                              (nios2_qsys_0_data_master_read),                                //                                                     .read
		.nios2_qsys_0_data_master_readdata                          (nios2_qsys_0_data_master_readdata),                            //                                                     .readdata
		.nios2_qsys_0_data_master_readdatavalid                     (nios2_qsys_0_data_master_readdatavalid),                       //                                                     .readdatavalid
		.nios2_qsys_0_data_master_write                             (nios2_qsys_0_data_master_write),                               //                                                     .write
		.nios2_qsys_0_data_master_writedata                         (nios2_qsys_0_data_master_writedata),                           //                                                     .writedata
		.nios2_qsys_0_data_master_debugaccess                       (nios2_qsys_0_data_master_debugaccess),                         //                                                     .debugaccess
		.nios2_qsys_0_instruction_master_address                    (nios2_qsys_0_instruction_master_address),                      //                      nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest                (nios2_qsys_0_instruction_master_waitrequest),                  //                                                     .waitrequest
		.nios2_qsys_0_instruction_master_read                       (nios2_qsys_0_instruction_master_read),                         //                                                     .read
		.nios2_qsys_0_instruction_master_readdata                   (nios2_qsys_0_instruction_master_readdata),                     //                                                     .readdata
		.nios2_qsys_0_instruction_master_readdatavalid              (nios2_qsys_0_instruction_master_readdatavalid),                //                                                     .readdatavalid
		.altpll_0_pll_slave_address                                 (mm_interconnect_0_altpll_0_pll_slave_address),                 //                                   altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                   (mm_interconnect_0_altpll_0_pll_slave_write),                   //                                                     .write
		.altpll_0_pll_slave_read                                    (mm_interconnect_0_altpll_0_pll_slave_read),                    //                                                     .read
		.altpll_0_pll_slave_readdata                                (mm_interconnect_0_altpll_0_pll_slave_readdata),                //                                                     .readdata
		.altpll_0_pll_slave_writedata                               (mm_interconnect_0_altpll_0_pll_slave_writedata),               //                                                     .writedata
		.ccb_slow_per_s0_address                                    (mm_interconnect_0_ccb_slow_per_s0_address),                    //                                      ccb_slow_per_s0.address
		.ccb_slow_per_s0_write                                      (mm_interconnect_0_ccb_slow_per_s0_write),                      //                                                     .write
		.ccb_slow_per_s0_read                                       (mm_interconnect_0_ccb_slow_per_s0_read),                       //                                                     .read
		.ccb_slow_per_s0_readdata                                   (mm_interconnect_0_ccb_slow_per_s0_readdata),                   //                                                     .readdata
		.ccb_slow_per_s0_writedata                                  (mm_interconnect_0_ccb_slow_per_s0_writedata),                  //                                                     .writedata
		.ccb_slow_per_s0_burstcount                                 (mm_interconnect_0_ccb_slow_per_s0_burstcount),                 //                                                     .burstcount
		.ccb_slow_per_s0_byteenable                                 (mm_interconnect_0_ccb_slow_per_s0_byteenable),                 //                                                     .byteenable
		.ccb_slow_per_s0_readdatavalid                              (mm_interconnect_0_ccb_slow_per_s0_readdatavalid),              //                                                     .readdatavalid
		.ccb_slow_per_s0_waitrequest                                (mm_interconnect_0_ccb_slow_per_s0_waitrequest),                //                                                     .waitrequest
		.ccb_slow_per_s0_debugaccess                                (mm_interconnect_0_ccb_slow_per_s0_debugaccess),                //                                                     .debugaccess
		.ccb_usb_s0_address                                         (mm_interconnect_0_ccb_usb_s0_address),                         //                                           ccb_usb_s0.address
		.ccb_usb_s0_write                                           (mm_interconnect_0_ccb_usb_s0_write),                           //                                                     .write
		.ccb_usb_s0_read                                            (mm_interconnect_0_ccb_usb_s0_read),                            //                                                     .read
		.ccb_usb_s0_readdata                                        (mm_interconnect_0_ccb_usb_s0_readdata),                        //                                                     .readdata
		.ccb_usb_s0_writedata                                       (mm_interconnect_0_ccb_usb_s0_writedata),                       //                                                     .writedata
		.ccb_usb_s0_burstcount                                      (mm_interconnect_0_ccb_usb_s0_burstcount),                      //                                                     .burstcount
		.ccb_usb_s0_byteenable                                      (mm_interconnect_0_ccb_usb_s0_byteenable),                      //                                                     .byteenable
		.ccb_usb_s0_readdatavalid                                   (mm_interconnect_0_ccb_usb_s0_readdatavalid),                   //                                                     .readdatavalid
		.ccb_usb_s0_waitrequest                                     (mm_interconnect_0_ccb_usb_s0_waitrequest),                     //                                                     .waitrequest
		.ccb_usb_s0_debugaccess                                     (mm_interconnect_0_ccb_usb_s0_debugaccess),                     //                                                     .debugaccess
		.dma_0_control_port_slave_address                           (mm_interconnect_0_dma_0_control_port_slave_address),           //                             dma_0_control_port_slave.address
		.dma_0_control_port_slave_write                             (mm_interconnect_0_dma_0_control_port_slave_write),             //                                                     .write
		.dma_0_control_port_slave_readdata                          (mm_interconnect_0_dma_0_control_port_slave_readdata),          //                                                     .readdata
		.dma_0_control_port_slave_writedata                         (mm_interconnect_0_dma_0_control_port_slave_writedata),         //                                                     .writedata
		.dma_0_control_port_slave_chipselect                        (mm_interconnect_0_dma_0_control_port_slave_chipselect),        //                                                     .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),      //                        jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),        //                                                     .write
		.jtag_uart_0_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),         //                                                     .read
		.jtag_uart_0_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),     //                                                     .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),    //                                                     .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                                     .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                                     .chipselect
		.nios2_qsys_0_jtag_debug_module_address                     (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //                       nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write                       (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                                     .write
		.nios2_qsys_0_jtag_debug_module_read                        (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                                     .read
		.nios2_qsys_0_jtag_debug_module_readdata                    (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                                     .readdata
		.nios2_qsys_0_jtag_debug_module_writedata                   (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                                     .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable                  (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                                     .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest                 (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                                     .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess                 (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                                     .debugaccess
		.onchip_memory_s1_address                                   (mm_interconnect_0_onchip_memory_s1_address),                   //                                     onchip_memory_s1.address
		.onchip_memory_s1_write                                     (mm_interconnect_0_onchip_memory_s1_write),                     //                                                     .write
		.onchip_memory_s1_readdata                                  (mm_interconnect_0_onchip_memory_s1_readdata),                  //                                                     .readdata
		.onchip_memory_s1_writedata                                 (mm_interconnect_0_onchip_memory_s1_writedata),                 //                                                     .writedata
		.onchip_memory_s1_byteenable                                (mm_interconnect_0_onchip_memory_s1_byteenable),                //                                                     .byteenable
		.onchip_memory_s1_chipselect                                (mm_interconnect_0_onchip_memory_s1_chipselect),                //                                                     .chipselect
		.onchip_memory_s1_clken                                     (mm_interconnect_0_onchip_memory_s1_clken),                     //                                                     .clken
		.onchip_memory_s2_address                                   (mm_interconnect_0_onchip_memory_s2_address),                   //                                     onchip_memory_s2.address
		.onchip_memory_s2_write                                     (mm_interconnect_0_onchip_memory_s2_write),                     //                                                     .write
		.onchip_memory_s2_readdata                                  (mm_interconnect_0_onchip_memory_s2_readdata),                  //                                                     .readdata
		.onchip_memory_s2_writedata                                 (mm_interconnect_0_onchip_memory_s2_writedata),                 //                                                     .writedata
		.onchip_memory_s2_byteenable                                (mm_interconnect_0_onchip_memory_s2_byteenable),                //                                                     .byteenable
		.onchip_memory_s2_chipselect                                (mm_interconnect_0_onchip_memory_s2_chipselect),                //                                                     .chipselect
		.onchip_memory_s2_clken                                     (mm_interconnect_0_onchip_memory_s2_clken)                      //                                                     .clken
	);

	usb20sr_refdes_mm_interconnect_1 mm_interconnect_1 (
		.u20_clk_out_clk_clk                             (u20_clk_out_clk),                                        //                           u20_clk_out_clk.clk
		.ccb_usb_m0_reset_reset_bridge_in_reset_reset    (rst_controller_003_reset_out_reset),                     //    ccb_usb_m0_reset_reset_bridge_in_reset.reset
		.usb20sr_clock_reset_reset_bridge_in_reset_reset (rst_controller_005_reset_out_reset),                     // usb20sr_clock_reset_reset_bridge_in_reset.reset
		.ccb_usb_m0_address                              (ccb_usb_m0_address),                                     //                                ccb_usb_m0.address
		.ccb_usb_m0_waitrequest                          (ccb_usb_m0_waitrequest),                                 //                                          .waitrequest
		.ccb_usb_m0_burstcount                           (ccb_usb_m0_burstcount),                                  //                                          .burstcount
		.ccb_usb_m0_byteenable                           (ccb_usb_m0_byteenable),                                  //                                          .byteenable
		.ccb_usb_m0_read                                 (ccb_usb_m0_read),                                        //                                          .read
		.ccb_usb_m0_readdata                             (ccb_usb_m0_readdata),                                    //                                          .readdata
		.ccb_usb_m0_readdatavalid                        (ccb_usb_m0_readdatavalid),                               //                                          .readdatavalid
		.ccb_usb_m0_write                                (ccb_usb_m0_write),                                       //                                          .write
		.ccb_usb_m0_writedata                            (ccb_usb_m0_writedata),                                   //                                          .writedata
		.ccb_usb_m0_debugaccess                          (ccb_usb_m0_debugaccess),                                 //                                          .debugaccess
		.usb20sr_avalon_slave_0_address                  (mm_interconnect_1_usb20sr_avalon_slave_0_address),       //                    usb20sr_avalon_slave_0.address
		.usb20sr_avalon_slave_0_write                    (mm_interconnect_1_usb20sr_avalon_slave_0_write),         //                                          .write
		.usb20sr_avalon_slave_0_read                     (mm_interconnect_1_usb20sr_avalon_slave_0_read),          //                                          .read
		.usb20sr_avalon_slave_0_readdata                 (mm_interconnect_1_usb20sr_avalon_slave_0_readdata),      //                                          .readdata
		.usb20sr_avalon_slave_0_writedata                (mm_interconnect_1_usb20sr_avalon_slave_0_writedata),     //                                          .writedata
		.usb20sr_avalon_slave_0_byteenable               (mm_interconnect_1_usb20sr_avalon_slave_0_byteenable),    //                                          .byteenable
		.usb20sr_avalon_slave_0_readdatavalid            (mm_interconnect_1_usb20sr_avalon_slave_0_readdatavalid), //                                          .readdatavalid
		.usb20sr_avalon_slave_0_waitrequest              (mm_interconnect_1_usb20sr_avalon_slave_0_waitrequest),   //                                          .waitrequest
		.usb20sr_avalon_slave_0_chipselect               (mm_interconnect_1_usb20sr_avalon_slave_0_chipselect)     //                                          .chipselect
	);

	usb20sr_refdes_mm_interconnect_2 mm_interconnect_2 (
		.altpll_0_c2_clk                                   (altpll_0_c2_clk),                          //                                 altpll_0_c2.clk
		.ccb_slow_per_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),       // ccb_slow_per_m0_reset_reset_bridge_in_reset.reset
		.ccb_slow_per_m0_address                           (ccb_slow_per_m0_address),                  //                             ccb_slow_per_m0.address
		.ccb_slow_per_m0_waitrequest                       (ccb_slow_per_m0_waitrequest),              //                                            .waitrequest
		.ccb_slow_per_m0_burstcount                        (ccb_slow_per_m0_burstcount),               //                                            .burstcount
		.ccb_slow_per_m0_byteenable                        (ccb_slow_per_m0_byteenable),               //                                            .byteenable
		.ccb_slow_per_m0_read                              (ccb_slow_per_m0_read),                     //                                            .read
		.ccb_slow_per_m0_readdata                          (ccb_slow_per_m0_readdata),                 //                                            .readdata
		.ccb_slow_per_m0_readdatavalid                     (ccb_slow_per_m0_readdatavalid),            //                                            .readdatavalid
		.ccb_slow_per_m0_write                             (ccb_slow_per_m0_write),                    //                                            .write
		.ccb_slow_per_m0_writedata                         (ccb_slow_per_m0_writedata),                //                                            .writedata
		.ccb_slow_per_m0_debugaccess                       (ccb_slow_per_m0_debugaccess),              //                                            .debugaccess
		.rst_pio_s1_address                                (mm_interconnect_2_rst_pio_s1_address),     //                                  rst_pio_s1.address
		.rst_pio_s1_write                                  (mm_interconnect_2_rst_pio_s1_write),       //                                            .write
		.rst_pio_s1_readdata                               (mm_interconnect_2_rst_pio_s1_readdata),    //                                            .readdata
		.rst_pio_s1_writedata                              (mm_interconnect_2_rst_pio_s1_writedata),   //                                            .writedata
		.rst_pio_s1_chipselect                             (mm_interconnect_2_rst_pio_s1_chipselect),  //                                            .chipselect
		.timer_0_s1_address                                (mm_interconnect_2_timer_0_s1_address),     //                                  timer_0_s1.address
		.timer_0_s1_write                                  (mm_interconnect_2_timer_0_s1_write),       //                                            .write
		.timer_0_s1_readdata                               (mm_interconnect_2_timer_0_s1_readdata),    //                                            .readdata
		.timer_0_s1_writedata                              (mm_interconnect_2_timer_0_s1_writedata),   //                                            .writedata
		.timer_0_s1_chipselect                             (mm_interconnect_2_timer_0_s1_chipselect),  //                                            .chipselect
		.user_led_s1_address                               (mm_interconnect_2_user_led_s1_address),    //                                 user_led_s1.address
		.user_led_s1_write                                 (mm_interconnect_2_user_led_s1_write),      //                                            .write
		.user_led_s1_readdata                              (mm_interconnect_2_user_led_s1_readdata),   //                                            .readdata
		.user_led_s1_writedata                             (mm_interconnect_2_user_led_s1_writedata),  //                                            .writedata
		.user_led_s1_chipselect                            (mm_interconnect_2_user_led_s1_chipselect)  //                                            .chipselect
	);

	usb20sr_refdes_irq_mapper irq_mapper (
		.clk           (altpll_0_c0_clk),                    //       clk.clk
		.reset         (rst_controller_004_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)              //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_0_c2_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (u20_clk_out_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c0_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_005_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (osc_clk_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (altpll_0_c2_clk),                    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (altpll_0_c0_clk),                        //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (u20_clk_out_clk),                    //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (altpll_0_c0_clk),                            //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_004_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (u20_clk_out_clk),                    //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
