��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��s������\�Ἡl-�y�f�����f� �ѕ:�nA�kb-q��_���ѹ(4�dê*���7��N2�ɐ��+ٞ�4Y6Mx�ejǴ�y9�����=���D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��\\�l�����r9s��@'�k~�{�<���y�#���i6`#Ɉh:^[����*`��Z��|���z���N?`q_���ר�Z���FLe���Et *�mk7���-��fP���� A��׾��o��Ӡlv�jj�����#�5!�����Ѿ������Rf��Ȏ�����ٺ�:G^7�A'�8�7��������J���А���W����i�k�d. �58+&s\9��]3z |xkbm�F�GɤD���zSl��x�za{����D2���5!���
_���c���E�;����C�6p�$8�mc	N����[$sq+C�o��:���vc9MR�|Z����;`+~�;"n�ԴQ@]\��R�|�4�ː�бÂ{R��O����)Z��k�&�O��7E�yM`>��5�m�"�^63�}�����8A��
+<�%��M�g)�G`:2�[c�Dw)x��y�'� �����m�v��DI����O鈩�0���R�5@��t��㒦�9��o!@& ����v�W���s��mnS��j5�Ѣ��lѓѱȦ��-H������t�	�&�k�M���4�!��X��#�x��V�p�$��ɠmsܓ
Y�A��\RS��H�
��}{s�~8�`��_b�f 1�a��9�E��pi����x|�&��A�8����:]B9/铪DpRqSxt��g˙��t�"*W�\���+��:�Ac�$��Lt����>k&kX���4>>:��+E�)%:���Dr��I������
h�7�U�-[?��Q�L���{� �,���12�(Йʌ��~k�J�����j������`�Ȧ�um�J,(l��ãM)�ׄ^���:PR��;`��2�@�i���7T��鄺5<��*,�q�H*ߎ�HR��I?��AK�t�[�N�d��R�l�v�1U{��X0Bx�g%��=d2ڜ�WLt�b%�r�-e�x�m��zlE�W������?��`ߘBl�	�vw�@�pnn��	%��;�PdGWO�Q3b7����� ����B'�Y�ډAy���&���E��ZX��	�u��UR��u�<m�����.�������dH�5�����[Bl�&�
S~Ch��՝�^"�p�����V<��.ӕkO�����
X����R�����`�����]�ݻ�M�HM
�X�6�i뢚52�2�J��@�cۡ�i�zU�4Eu8�S�� ]�o�������b׋Ao@��ѵ�>� �"#���ǽFe�����e&���$��r2��x���)oxV]Ȅs�"��1!|<�Ͽ�iE����D�V�p}>�4��P/�"ʮ@���N�$eM-DRʌ�)8!�"�ҖRPH����QB�AY�������9I�Hq��Gbղ�ہVl�4��RV`�׭��-�X�S��6���T�$*^�w"�X'�!�ZwFl)z3�X�@*d	yM%w嗂�٪�I���$��v`�5��gSb���� �T���`P��0���B���ה��]V���fa�=�l�s��{��	���:Ε\}������Ro����DQ\�uP�%;�̏��Ta0r)$QVݣ1���N��M{���*~a�ybF�kZ�p�vb�:E����x�(�ţ�L7�����O0K���s�g)�3cV1�L��q�!��Ӽ4�i-�N*n�/i$6M�������f��)ѩ\d�)�5;z���۝��x]Z[��p�+��U�>=�Kuq�a�I�3	�U�y�5u�k�Ѽ���{�����f�|�$C�� �~� 3�U��×a���fgO	��	����m���A	�(p�J���l����j�/t��R4�x�?�k�1�G]��h�7��&x\5�˩|`����~�Ւy6@b�n�k�.]�������P�?)�7ho2y�&��� �	��m�b<&��2T��^Dgc��}�5X�y��|.af�eA@�qŊr��5��Yw�]���_�5��Er��>@t�RC"+9P��r��q�7��le�\��8	�e-����P&�o?�}i^(�V�#P[�O��Ѱi��y�t����Q�ǟG��� �_��T:R�S�/C��s[��d������θ��`j���s��L���̬�y �Ϳ�9��*��W��/5j�y;3rKHm;����Z��$�H����DJ�$�,P�J�F%&�ۖhƫ4¾3����|kx2�����LQ�Z�W�T��v~�0�!�C�������07ס�TyW��iR��J M�A^��I��k�B����p�)������9������`y5���9 �ـ2�gd�R-�^�^Η��:�sG<hv��p�a�Ļ�,隸inN�ExOp�	v�M[XE�ޱ3�?.��! A ЭG���wVFޘ����BN7���Ń�d����fTr���p^B�j�N���Z���q:��ٜǣ �!�|���_�ϴ3�}��`F��Sz&�#�m�^
�S �Zu]'I�c���ɔ�d$9�AN�����Z\L6��A0��K'IX�H�O� ʲ�Cj�	�B���ۄ�ǎ\��(H"^A0`ل��46��Q]����b�)���7���f����Z��@:�*˚�� ���xM�T�b�~�ll�P͘Fs����>�%W[�@Ja�!C/c� �Ŝ�F�,�R#B�BΔ��Y��ۧ�T ��1�,ɩK�1o,��}F�u?���Zk)R��ˋ��+�ÅW�-�"��g�����Ȩ�}�?��Z�㩪!?����o���E�Q0���2�'�W�!�f�����I.�Rc���g���e�4�e���%j3�{���g]6�ޮ��$p�� �)�x4�Dv#x^�X<��Q��y&`�J��!"�lJ�@+��b3{�h�E�d��R�9�"'�r}&���Qnz�ݡ�J��5��>�bͤ@h��P�%ÿ_7���@`�P�҆N���k�����U�6j�O�`�g?$fԭF�M�_�dVP��m����������~^ne�A��eg��0�9Q8Hs곬ZW�g�T��Lf���P���pL�
K��Y?|��峳�}3�y����,B��� Y�����:�}�d=n��	��PcU�8��(��%�|#_F=ORZ�%�iS�����'���K�Lvt��b��c.%���]0̷�Y�]
CҞ���M�േ �Vf���1�"
�hv��O0�gҗc�5�]k)�N!c�W���#���q!�J��3��ݔ�5�2KW[�2[ئ7qj��!�J��\%��KĦ ��K6�yM�;�r+[S���e��{��p�Ĭ�h���r�X�=&tr�]��!���%��?p~^�����_8������\op��v�B�b�H�l5���ZY� 0���� A%��Y�@������ΰj?6���Z�bd����Hu�@��"<
���P��˥���kx!�c=���]�}�������d2�moږ�iV3��<����$.���'f��ꧯ��Á���msA/>��;�� �u��tB�^�M��hq�ڮ�o��x(92Ia-\��=�g�g�
�E,9Q�Lֳ�p't�͸Y�b8��{�+�ͦ�{��ۦ g;�(�����+!��N�4Cz� ���򛙣�� ������^96Gxڤ(�a�D�7���o�����r�$F����w�&|�nM�����6�[��1���.�p�ϳժ���1^��Ѓ�T쎫���v�N�x)?���Q��ء��y���>��p4O8�/~�������}�A�X�%������i����˺���/&�Y�
�J�)BT�g��EYd��@Ho�\|�ˆF�7ࢩ��L�>w�^�LG�-�
���P�9$C`��/oU�y�6��<��KU�f���`>c!�?��#h"���������S}�w5������Hc�4�ݍ�9dwm���}C4T�'��a�����|��t����&�d
bb�鞺zcP��N�bјL����5^~%V�]�bY�`�-*�:c�|�K�#�Z�g#����ra�~�,~���R{��e���tR�s=�;�K��x�y�ؼ��v����@�|�HN��׉z�_��������H�&a:����3�P�fa�'��Z��)kU�\��1���[f�e����6�i�"��2�|�~�C[=s4�f��f<�T����b]f&�]Qq� d_Bٴ\̤"EN�
:Lm{5[�������ض�v��[r��=�G����� ��襵�i�;ůk�@��и��֕h=��4r�_�����kB<���z��21d9Y�-��-��~��y����u=	D�s�5\\N�k���
) ��5?A�e��O?3��/�'�O�Ɲ�,�6^���WUh.�װ,�����Xd�^�7N��gބ�!�o�I�!>�K���D�Br�S�<�'0>�m��8��dwi��"S�:[����q��ңpR�����֕G�q~(>\�,�O���\�K<V&�v�k�V��?��$�dP�,@Z��h��T׭���n9�bn�����a�y�	*J�9��n�0�����"��JsP���D��)��=-�0���ygzyЍIt*�L��h��9�<T��|���K�n��g�PԺ�T�m����7og�\zG�(��'1�����W���KQ8_�o����Q�KT�tDp�_T��E얂ډ�-`~�* AFPu�]��:���7cL��A���ka8v�f0%�6"4��j��ܟ�M ��c��&>~O&՝�`����sTa_X�ŝ����K��c����H�B��p�AzTK֟��!o�*HY�KM8Vr�̯~۬����rܙ�o�}`���?� d�����-6���o�!u�:?��&���f_~�c�<{���&�hs� j��H�5���.��ɱ-*G��n1�%iH�����"��^c�y���,
������*�Lַٛ���qv̪�%Q�~�R�J>	��Il���=��jWܣ���`Ʉ��C���b���Nr�TAS��.��v*�Ppl�f��lǞ�3�5��``��B�hr�v�3UlN�A���UT��{Tyk�@  f�l��S�M:ڜ��yT�]�afc�t?��`,m���h��-* �&rO�h\��P��:����t���D-p��)�_�(l���6>l�y�̛��U޼�nt2�0���>T�Ni�ܣ�$1w�w,�=�u��E�x��<b�o_�|�, K!��B5�	�9����7*5�V}b:�e�%�5�7�@�����ܝ�K��4��_,g��ٜn,�����rXn%�(��ho	e��ۡ� �t g�޿8�C;p��j��d�Osg)d�a�մ�%��V� S7O	�.�37>[�a����N�X����.X�l�{���u�c�E��<���uӬh�:\]2GȨO��7���r�$�C��F9�,]���j�O���Q��\^��S��mnϮ����˩�e�QS\�PR���5��d�>T�X��aT?Սz�j#�0��k�l��XAg�8�^乤�6q{O�������ptƭ�rf�>#�ԢI�/�s�P���q	k�J '\vr�%~8p���N�����'��u�de7� ��/���$rc�0���{%╩��G��خ�(�hA����!v�Y �x���]~�,0�HD��X�\����3Cet���tln�ॳ��kAIrmG���]�7Z��b�����w�*��P���I�0��k�Km1���I��굲%��bM=���ǀ�|:�r���%lK���	�E~��#A��[׿�z�[�;��z��zަ�w	y���E�:W�wH@� e �j�2��+`u�;#ԕ�+D��_%/�k㐥�\��Nx��c��b��t���)P�u���sl����lSj���w�:��U�z3�(&���2���0!^授������Zx��d���`�9�x� (�B �3����p) x���f����̧a���o�&F�����z��vp��vҜ��^>�~�]�=�($u��s�NY�K���|�TJO�`B�a-�މB6��2a6QSb7�`��[1���� x4�� "9��t���,�VQd��N�z��p�;�f� ��.a���>آ(�|#YC<8�'��� X�7P�+�x�G�*�)/4�l"?������#��
�XP�F��C򦝋_��A�-E!͙h��~(kȟ��*U1��ϼ�mP�I�
���JEj�G��=�-���rڅ�{:���Òowm?������V^�����p�r�9
�}�E��LqCG�j��P�<�ލB\� -���QkIW��6���~L[��x��i_^�P&d��Y�F3v.�����Z���u���P������e�Imc���4C��k���f氎 kf]5j�3��ro=�;�����]|9�����01���G��c�Pe��4��>S��?��{�E���wNDg��u:�����$\���X{Xs�`䉫�p�NE��Z�*��w�q"خ���hI~�H���� ������O��M`͛�Qo|��E;myK��Q�3�����LK��@�|��Nj4�B~��~j�M$���ƛߊ�p��Z�g�A��1l���2���*w��y]�q�B��䟒@�	d��L�k��:+\9%�眬u���m���Ї	�`�d2p^W$�P[A{�P�;]x��#zf_B���ut셑��kxF���������E|Ax�K{i��*�eoy��]5�P2o�M�>-��D��h�W�q=�;:����!���<H�m��i���>�Ϸ�ĂX�� ����AG�>f������3�L#R���F]��6�&����N� fMVR��=I�<�qIB�Vf�6��aL��=s{0h���3:|���2�?3�F���,�8%v�P��VK��O 
��Q���֗3�$y�<f�2R�Zȣ���AYD�C�K�v 6�2��`�ܠ(s+'�$zѫ���J,Ou���ɘ8 ���W��Sf%[��=���%Xdv�6�;�T�g��G�H>�cc�-2��)PxR]�fvP�r������@�P��誹��6+��\#a��z=���z��y��w���h/f��h$;z����Tx�o��45@0��G��/5
��P̮��$�����Q	c+��e�Ń
Ѿ�N�u\2���9�9�;x��G�(� ��`���Y����3��KϮ�0��ʫ��Q��Zk�l+�\�۴�&B�A���	0�ʆ�l�"»�F$���;�pW���0qB ��D�1&�(M���"�����705F1ɷ*jeo���XȪ�n�ce٧��͝�m��dѺZ/��#tu�O
]�7�mIN�N��L�;�<�C��n�qV�yʑ�+��e��� �JÞg{ir�p!1�ÿ�;=|��V48&4�O	��X�R�O�[��$4�V�Z�h�k�̭?�
����NUz������0���ײ|ѥ8Z�S\��7 ��t��)J��M&9q-�RU�v��歈�/��%h�'�L�(�~�"��!�3��9�F�D�E=3a�v`��r�{Gu�4C����:ך�h��7
� ��햗3���<�����GY�)��nk�ϴ�A��Cyw@Qz��� �Ĝb��6_܃�ɵ|΍^�7d���]�������5
���M�S��!�B�/���h�~)�t3�i�����%z:E����,��/�XN~Jp�פ���K�Z�Q���-_
���j���A��7���'��U�	~,��h�2q��D
�{�dB��,�ؒn�et�=붕��
#��ܲ8��y_�%uGtņa����.�A������X{�X"N��:��'R��H�_��[�^��	s��=F/YCtC�:4����4�r�"&hP�'�[��nzn���E�e�
���:ټ��p�SdE���dt�a��x�\�k-�fJZMX	�B�g�"Bu�M
�Ȼ��t����@>�����5(�$* ݦ�����_=ֶ@���UҨ�E��n���S�&�����p�-+丮M�w#�N�&���$�B���+ �<0�x7_��> 2��t��(D����\�/"[X���]��C��Ct�Mi��=a/U�WA"7�w|���M��V����9�t����wQh#��K{�A���)3��}�y;��X��W�D"=�����p���f2`���z���Vc�G0�(���J"�.<���p�����ۦ�髵T@�ޯ�z4��bv�{�qӞ�%eD��'�~t���:IU�A�F�$�Q�x�����JT-)AѸ)m7�����!}����#���nzB�j�]�w���[����0�*8�p����Z�����-u���-{>of�X����D���0�CK˲� ����R��y�p�G���b��Z���
�I�'�������
&��ۯ$��W�1ܲ�k�=�P>�U5H�]��P�NȮV��9ӕD��s�F�sd%W����ZI��Mj�����04�J�(���� w����8�Rq���8�tN�K�C's��'`�{ţ6���CS���&�1�$6�]6�^��e~����0*���a�8�g�zߢ��:����2�;{v�l�g��)&�2dpXH��]c�T][)�x��ȴ��)�b�d����'h���yN�a��s��O�C$�'��ރ~4�TL;�YX9%/�o��X��`Ά�~�:Շ=�F�����7�H[��\d.֌j4g���#!DV�-�*_����1SU��{y��7*
c��9�J�9m���B�1��j��"L�!Aˀ�$!�?2���̇^u"(q�^�9c��g�%������,}V�g"���rq�|EXw	��q��T�z���uτ/����LǄ�$Lh��K��k��Q�N;|�Ԅc���e�)����~�m�@da"�����9t�\}�n�˟C ��L�f"� '�DgN]L�3�FK��Z�g/Vc�+we0h��;��ۃ��'Q��:i4M|J��P(���ɧ~=ݎyG��{ɀ@�D�_�?����.�Êg�{��<�Q�Z9SH�����/9 �o���Q',�%�[���<7�l3�)n�#H����%_��z���ӝ�3�Lt���nLll�F���3��:"	�s-3�H��%k'<F��'z2�����*j��m����扊��|ǟeh��� �p�*x��n���1�(��V$,�lv%ET�p���Ē�τ�B`��^��a�$�uJ3��]E��F\���P/<��E ;}[W�Q�fg����Fҽ�]�Yݵ��{#{r�?���}�:�
5��&oB�0V�T�Š r	D0�[\���&��m�*���5�_�_�m��=��v_D�B�(4��cȹ�6�����r�+n�Q��j(����`O&��X����E��D�R�"zV��)=�T��	v��-�i�֥�N[�J�u�R�Y:+6h�K�jt���C2��~{� ������_(;��I2�is�6�9Є���^D� pο�eq`��Vו:����乇Z����"���g!^�����1Uj.�~�$�h	��ayz������f�h�)��93ǰ�S���?P��Y �J��|�#���Do�(,���t�vW�&�������s�rta���Ǫ;����O�{���G7z,�yun�$���BӅ/�=�Vzr����&t�Κ�4t�u�Ώ�c�9�X,Bun�\+����F�c�/e5��2f��&���>E���������KF��<�gDc�k��3�wB��������\�6�s娎;�Jc 	w>6�@Z�xr5��gə0�#�=��*�� XQ�P%���ujr3*a���j������4>B*;��4
�0W7Kk�A�@])�����Lz&γ�h5r�|V���;��*���	MQ7x֫� LU�t/!�j�� J��N�"IJ�����C��B_���|�:_��BZ�S�^D�q��:&Y:�-J�a|7�YȹZ#4�~W����"��2<j��4MT@�?��n�0==K�G��_�v����#��/��$���x5ߘ�}���pG|v�y��+u�B��8�m�L-Dsc���ó1]r]�SYW���*�s��f<��P�:�Ԋ�B3MB��}���7�}�����?cj6G�BA�6���"�-Ԗ��sr���KwCn�"�3�Q�a/0�
ռLJ��``~��%$�k�6+��.���kYC� ���N�	�h)��8�㫥�w�R64��7���ȍe���'��٩��-\\V.ť$+&f�X��c�绞��"Ä�X������"]S��1c�y���b8�ˈ����)T�C �Cp{(�����WSؿO�)����|���D���`�����Tp�N����+7�z����}��l�U�ò����˺D�
3"�]jk<]^����lw�®��(�s}�����hG�e�4w 3a�&�mտ��|ڒ�M�;��"E3 M��MjK{��L��� 	aK]x�*�>u���*T�l��2��U��ٖA�#���L��	gO�8.�A5�
�
�;��4@˶�2�LڦXoƼ��پϚ�~���R�9�;�>IJ�\�k� ����0�M�����g��g^�j2�fRWb�~��@e��'`J��M G=U��/[v�
��n����$��R�bӈ�ͩ?l!��Gzx���2�](��П����= 
B띲&�Z�a��r�xR,#�Ln�Ӎ|���y?��L���������ڃ�����5���O� v�VӊA�Hfu�
�&Aݜ�Y�Y�(%e��;Ι�e�T26a�D�>����R~19�BwI��b�"�E"�0�%V\�-��~�W���*v�����H�Hi����XR}���R}�f�h�Xj▸��'�Lg�"�||���6b�������|}8�;&s�-��ܫR�,� [�:2$��Iꃏq{�	+��_B�K6�3�CY��~f����e:��B��*��\c`���k��E���0��֯*=�{�aӕ��"�\5�\��P/ހ� 3wp��x�����L��^F��"��C�P%3���0Q��w{�1cEf�W�/���w�Gi�=K�������U�c>�{]�����ˡrE~6gt�#YD!9I���O�������������^�/�AU/d�o1�H�Bxn���_�A��p_�{�ˢ�1Ym��Rd��@>b�H&�.?+è�Ӏ�y�~� -SJ������h����W���. i�A�T�Sa.8���K�i̽\�W�L0I���~��H�X��$|+��e�($��l��?��g�JmVT�Vt󾜼�v_!��x�{f�2T���É{���o���χ.,����3�3?�)��J��&���8cZ����sjZv�lf��� ���2���ҍ������K�2e%2����gX�ϴ�v��ӹ�T������m1��)	Ҥ��=�IǞ��޼�G��+ ɥ9U.K.$�����`؇�ύsN�q�%��uy4�jװ���7y���4u�,y�DsSU���tAXg::�9<G���D;c�޹8Q��z���	:���m���b$O{�|���r�\�sS5�
T���܊�3��|Sh3��5a!��6�u�|�ۼ���=={}#\}���^���3�����:���q_�D�ڿw���z���H��h�8yWwG����绚dK�(��6��`ǒN��� =^����/r�-W#���hZ<1jl ��s�=� �(��K'�#������د���w!�������q���F����%c1Z�D�>U`L���k����yn�Ʉ,�vt��|�k�ʐѨ1����^���Ɖ��b%��=�/��{s��jNg �V{��SV�&ĸZ��~�66���U^`��L��]�1�vY3�������\�B^y<�R�4��r
d����8�@D_��XN�k�%�-U� K'�T8+��&G�0s���+]q������w"���Ό��w��S���0'�A.���06<��ƻ����_Q'z�2N�� ���noG��b�^a�|J3P��]'4��� �{�³���j,���L|*Ŗ{��[��a%Ϣ���m����U��h���Q���48A��Z`l3Rvi#�p������t���e��/��F�-Bo�6SX����"��X��Hڶ'�$����H$�[����z^�=��,h<zO���E����	���OӴ��y��bL� ���s�Y��gm��F�*���C�0��EX�ue�c��h\�K3q�ш��V�xt�e�@Y�5n��#��s���}��� kyᦅ��?%�������hh�|�q��C���$[y}N��~�qϒ��T�۹�Σ��G����u����_���8Rꅾ�Db9`�>e5�T��T=� ��9Ef�R,b�&1���[�9�T:'*�֥x�\'N��EÚ�}hw"��ϓ�1$Q7�z{�и��/G����[�BP ҂�Qpf��(֘{���Dꙹ��g��,_��9��#�w�VI?\卫Z�ygŝm��u5��9�&�� ��$а��JMc؞����.�ژf�3Ѹ�;u�#?�^#&u�����̪��&[�e�>�6�D��W����B�|ak��N����g�!�bՆ�)��s8V����`��V8`����s�^�~d;�b8����p�?`oZa� 4ޢ]�#o+w}�^@�D�Ic�3��Y��Ca�M��^�O�`���3��8��&I��e�5y���T,�	���t% � ���A�=L�H���&����a��O���~�)qs�]���:�0/R[2��x6����Ga�"�i�Ou#is�wS��:��#-�R.q��#��4��"I2U�����e2f�Q\��}�8���}��	I��x�m���M�E{zn$x�˽����UG0��q���D�l��"Z������d_��m}�2�9���Pz�j]`Jn~�uu���*:�Ԣ�ƞ�bV�����^��nK��X(�1���m�0n�y؏k�;�y���\7E̠Yi�&�R���{XU��U��Zyc3�aD�,��V�W#pO�����V܋�}�a&P����$�q�]�S��o�J��O"ʠ���E1��{�N�f�;��������-P*��z�ҹ�C�5�K _bF�.����KM��Lɋ�?P4��-u�Ge�g�Y��08Z�HM���>���%��e��[�>lnM�6jҟ!1��6u���v�-HK��>�}3�0k����A�=yq�Ǫ� �W�׃�^a�ԇŁ�DFs1�1�p�Rܠ�A��q��ބr�?�	>'��g�([R�!�&����K.){�S!Ȉ{Ad�g����ֻ��0�p7Q��[+�[j�v7!��%>ED�;�(q|N[���
���PT�y/�r4� H}�h3ł���CL/Ik-YD��!��-io�Q��k��G�B	��~{α���^<qM�H�+�z����i3~ӸP��B
�u��#v�5y���\g�5"�G"�\o�ks�A0��i-'���{n#��Tjx�g���߇��5t�W*N�G"C�c�)�{����$_[c�¯̑��U�]1�_�@Aƙ"��7v��݇�(�?B]*\24%n�؎��x��M����qIb������|�T�#ʐ\Z��?w4���\��˨N%~#0�B�҆j�8,-gDBNb�_Dy2z�v\��y� ��1s-�+]�K��I�w�6�x HLfa�ɊQ�c֚�JT��bf1׭�P߉6�U�x8kǶ��4$U��F"0�I���]{hoR�r*���b5�ի6	N��Ht��Z����_0W����ݓ���3��<��q�BO�C����������Rٕ]e�<Fo��!�敇h���~R89����	J�p�W5�Ο�3�զI>���^�L��_#U�������6���M���]N�~�et��/A�?=9��`Kh�ɾ񺡠X��]�)&U��|u�d�
3������p����_����G�O�篘��B�}�fb��T}�*��M�a{�����\]\�'�4�+]ţ�W�����o|'m�T�(L���*L�%?�����k��7|�EZ�Эu�U�Ql�]�:����e_�~E�ʃ"P	�a}��V��m�X\�_�=RhpĮ�?k��f��A�L�N3��,�w�.�?
�^��R�'{u�̘-�8!��t�,�J(�a�q�/b�w�\�z�s���y�/;+�N펌L�X`un�T���(����Cj�M���"Y.Qq���Iv�z�G�|I~�r/?�`������8�+���k�u_�����ɝ�A�������_]@�p��w���F�G�����$u)0̏�J �qio�f(����^ޞ���a��rP�p �EuP܇
'�p�=ԒdGR����A��ZNn e��^)�frf��i�����!�@Q�u�ͤ啫������S�y��V�%璣���$����~�J�(�5��@���Ө�7�EǞu=��jfT'�	d7ԹY�&/���I�+�F� �����;�i������pQM%/#:qn1E����ޔxz�I���Ļe3xG��	��["�|�b�i�ꅃ�=���"r����Qd�,i��`@ڒ��w�6Xb�^��'P؍B������
o7��z��sK@Ǯ�:���I��簸-��[������H�sUA�/��e�#�& LQ�2��1�!қ;�|A�&�PD ��0e��v �6���x��ys4����"�$G7'1#/�H;y!�"��x3���Ԟ''�Y�2^]���1��ӌ���0@�,}mI0G��y=E_������(0���ɇ~�g�r+�5�I��*A�ND
a��ԏ'0Y/ډ�Z��]�7,'B�'A����h�������A|���6R˂`VWU��&n^��`1�*or~��
9�e�e�%��p�U�5W��6j�������ɭ��XJF�Ã�
�1�%�	3��ꗽJ��������)��b��=�-���c�_��;�]��+)$�UkiN�Vq�QD�S�p��Ǚ�Ɩ_s��������ۂ��;���Q!��=_��u�К�p57q����QP�O��N��EH�/UN?����.��5>�6n�(�2i�W�&���v9��P�	Qg
B��(���e�H4i��}/"���bⒶ20���ل~V�ш&+�\F����Z|&V�쇮�D!]"6~na&�MB��K`{UO�i!��^@QMtW��XŀT$)�$ՒF{��������f���rx��ѢE&��#� @�}�6�߃I��J52HL?R����_�����Ḋ����������60��hgR|R2�<�nR�`�PT.��AHV̯5B���4?�k�-����p��� 2�-�߆oa���s�����8f��(N�yӏ���#�Q�Z���ӑ6wl�M�N�ZMW�i�U8�Y+/V�f.J���LA6�6&�Ų�/yo�k�^�5͍eI�.�V�W�-�ʫ�o�\x�/�Wv�a���ҽ���i~�a�o�,;q����bf���;��F�?���|�U*h��S�?S�+>��{�U�G<��\��)d��!��Y˝�{D�hOP���q0����o7��Q5ENg:��P�Z4��ΒQ�Z��v�X���� ���y@�^-q�U�T�J�P�����&��Ǉ�(�΄�e�ED�~_�@&0>M�Q%���+"#��O/ȡ�����2ߍ0�Lo����^&�d����9b=��mZ�^���q�ʑd0��U���bS����M��U�)^1��-I��ގh���/G���N|jo��'Ri�i�%�ea4�7O��i��-k��)��8'�)<�/�Q�f�A���9� ��G��+�DԱ�=��$v�7��u;���V�R�!��yۭUo�0� r	��i�Md5�2�Q)�o,#p�F�긴�B���1A�EE�\�z�����g[E�"%���Ad"D�B�.P��x�-�����3���0Ќ�_n���q��͋����y��%7�,Vg2�����~�&Z�~�[�]Q���H���T���J���t�W�A�"���d�m�.���ig1b��JYn�#G���	I����ls��[`���uy�������\a�p��C�u(p���&��H76����b�X{�l�&��S���t���{@+���3˪@�ܥ��[/{U*>}T��l�w���9��@<��<��l,���9����Ţ��푱�������wI
��VJ,��R���ZK�rF:bK�q)����̾]�fę�|}��wd<D���V���
��?&f�Z���Gcz�XW.��pݽ����hn:��K�n2����ݩH�l���&���n������
=��}�">xIV7r��i�nPC�Pr�������W�YC|K���_����������bω�q�#Cf�ʣ��2�`���@t(�p�:�LG����s&�&�{�ABlD��Il�g�~�K8���2jH���ز\��I�oI,���yi����ѷ���#;إ�=]��$tl+L�1����zHG��(,�5�p��	S����yF���eY[PmU�!�������鉔Ť��~�]j�/+��ܻ�{1���o�	���PEN �-}0R�b��˨���&��{�����/BYϩ��(HdC��}���r����6���p;V.�Q(]��Y��L#��ův@��YӃ�2�XW,�]�<����"��ޯ����TS�����b��
�����a�>(�fq#d	)��Jd�nV+E�)FK?�DD���꿄}�_�����Cp�3��۝�����q�3�����?[��
�+.��)�������+���(�S��T�4��
�Ս�iV��7\��z(MP�9�����9���F��Zk"�q��p&:�}a�Jy|{��S؊��zQ�����0u3ld������sX;}ْ���	��T�?b�6����Y���%���h�M%`����p�y�Ն�;
ݘD�b�2������(�7G:\wS|�Ylt$jU볡��:�˺�e(��&�-�J
k�u8h\b�҇�+%|��'t�t�ڼ��l�hB�Cl,�~C�7`�˄r�?���<� w�����%����MO?0��	���%˙���R��` ~��b�h>�j�6mm��*���[��:xUԛ��"1��(@!A�Ă���d�#$-�/�X��G����S��{��;���������E�1|�;������GR�L���-SL�O_��"&���E�-2��T�+ΐ��.�NPM,�)�]RփzA��v~��7��/޻!��]�iG���$�Q�KMb�{՞�U�˸�Y�ݩ*���
��T2�ǚ�o�NH�g]!�A�>g��g���5cGK��iO��^8�k	�+	Q;_J�v�ϖg�k=OĄ��j��3B�`KX�Y|t�vO�Z�� �։�(�R�=�8t�)��W�J:�)���w)5�R�.�_B�K��Q�ϛexv1���:<�׽�o�pbPN/��v����m}�����ߨ��X�-"~��R^�Nz����͝(Z.����&tO��IJD�Hծ���Ãk�ȝ1<p(z�1l����̪��Kb���2B�N��{o��茅�������#��~��L��58�z�ٚ�y,6��'�m�d�p)x!Z����:��]J&LPH�1Գ����>?<x誚"J��_�9�_`��S϶�m���QT;4�o�z��$=M�ϭ\l@�"���0�r�F�X��Ϧ�yu�/{�$;��!!��H%8Oڜ�Ϭ�K4^
7�!�3�(3��l�g�z�&۱���I�?�,��Zi\e�Z�/�$��%�өd�D8)�I��$��-z�ԥS��-���q�d��L%3YS���g;F�$�ݔ�ڣ5
;'a�,�|}<�9"��$sWbp� ��0h;���	�w����t�E���">%��?��
 <v�%�,3.���Q�KI�f�ës|����H`���z�h��mJD/eŗ$��݀���_��J^X�Y�>*'�xy��/#�H]خoRс�2Op�Zpy�{��yY�K�`�ZL�8π��2n���[�ry,z꺧�YmV�����!������*�5��	���Q��S�ߧ����pXQ���@S�Sl$��g��9����	{-�IʏX?ϫ���$H}���я�ECS�}��S*7;��֯�if\(�6���OO�$�a��Sٛ&�a9@F R^szI1�J�2�Z�9?nm�{���Px�}NPguD*�%P���W2)~*�{�����cY�t�*�x��������nfV@����!��4��{0(�:$\Rt�E��Z�'�OI�v��S�l�"�e I��?W�;���O�{=졒�9��M��c|i�����{�����ű��s�ޡ�����\�JK"pB��C���������_�u��-�e���V���C�g�0�8Q��m�xn���깎.M���7�H�;����CR=q���͎o����7�� Է�t����h�cƌ��46�1�7��� �D��S��厁F���@�����ܿ�G^00բ!�	}G�v��1�� M�n�`(`3�8�:#�oq�1b�|W�s?�M���s���8J��u�}ʵپE�2 U1Bkay��b�P	�|�|��������I����/J�Z�՚�A(!���c��
�*�G���ʬ"N�u�*�(_d6@4v�BY�*,\����	� Dc4��_lu�������C٥٪u�e�S���f���U`��;+*�}_Ϗ�DYG�~�jnS��Ɔ��v����Km�nI�UA��4"o�1�W�yz���%�ҥ�|�)u,l��k.IS���>�i�]G�D��O���������L}�������_�-��7l� ����w\�z�,�,�U���y).��@T�� �%�&���P��yֿϝ�B<�8������pnn��)s�� ㋧uM|2�Aㅆ����d�E����m3<:&/��5����~�eQ�'h��s�`Ι@1�[t*�2I����P*��4-��$F�MO6��x� jٹ���^��Ҝ2�j���{�����e ;`��h���H}��"b�"2֌X���������W>�b�'/���"v��辳�_|6J�� wC��(+��#���$�whU�(p	��'M�/�(�s�!ɧ1j
�C��(ƍ���SM�H���M!~F����p�b�̗����l�5U�oX�h��ށyv�+'t׊��[�.l��|��B�.Hse�C�G�b9Ǆ:�i��pw䣰�@�O1g�O�*W�9V�����C�����ј�;�����h<1�wŘ����P�� v�yK�ŘX��(�\#Qy)]�v.���w ���P+e'�}=�`����<��_	�|A�lQ4$�����0X2����� k�g�� �,���i�wҠ͢� 74p�b�7|�~��g��y?�I��}�9%���>����F��)ԅ]�|��Zx��c6��"�dVF,窙�kc~���V�̣�a�v�okM�<ij���&�i�Ȇ���z4���ޯ�����e���<c��a 0�ƽ���;�އ�O��x���6���`�G'�Ψ���� �9�U2`҅ � 7�)rE$y��\�j�s�r�@e����	�jj��x[sF��+]��>�A6�W�K�����aݥ��=k��;e ����J<���ąb�!�Pb�C5��#UO�W���$�K�>���Z�s��=x`nV|*����o�W�7�}��4�V��GC��}D�$E��Z����wsΡ+;�1���-�|��<wg
���^��I�]7����@:i�sv� �&DĠ���&tW4��nڤ�f@kZ՝z���`��]�(jA\k�z���ַ��k+�K�.>��&E�T�E�L&����J�F�^weX;��wu�,m�j_Eu�.�H����'���`W��Nk�#�=�,7?�:��ԕh���QV�x񇟝ԥ��<X�a/O�L����ր�9�Akv��@��ߪ�Rx�{v�w�E'�g��L��+vFL���J�"J�\]�w���и�۔G�6I��@�nD)J��K�Ծ�w�s� �!��:���B�uEd������0���(��}B�����m3�L)���\�V��G�Y���lﶪq��� T�)����y�������s�M.aΪ;IT�6_b������S�n���u�������u
8\��D��@Դ�#��4�/	��&d ���2lZ*i�>ta��e���[�dRz؛4Pijm,��z� ]�FI����o�;���}=c�YcY�id���?>�	>.Ԣ���;A*��v�ҲL� ��Ϗ�ӣ��]�L�a<4
�3g��m�����i�FF�$/��V|
��zُ^����蘤�+�hY�܎?��l�]9B�N�-%�
�#�߽�F�1_�V��J��l����D)����S��>م����MHU���eE�륁��u�/)p��`+�>y��!�����,�:;#r����=C4y@����hU_�42�!�:���ę�v[��� }�6UtJ��u��x2ز�����=��{q�b�C<&0�ɓk&��QS��c<�M����?,;�F[*�j�Ч�!M�@]�[qQm�j�֓��z<=����~�'�o��ed�m�Щ���v�V�SZ��6�f5!���y�zq)�nكv�*fl�@���ړk�g3�zu.%iq�,CN[��o+Y�XI��rϙֶ�lvN�@����؏��������4y�3�*���F)�o�'�x/>�h$��'�ݙ���uT(�bB�h�!L,K���S��Bk�N[��.��Z�7�k-M�+� 
� �m��w�=�{)'H���>��[����+�����������_�T	`ꂼ(�������F^�����= ƨ+�^ �aQ�W���5�.u�r������g���_��b�)�6[�)�F���"��q����*L1F]��G��w	���e���8�Xs��@pK��2��,/�仹�z�`����\t�w�i�3���������ـ̔ʥۙ�UvA\Ӛ5��3Z������Bs�.�;���~#hN��vj�uZ�H4�l_�����q��&a� �<�؜q�EM��BmK���5�^�,�5�,@��3��̱�OX$v� ��-D��,gLnxQ/�g�U�J�ڳ�I���s�k1X����ʄr^A��J�L��f4�7�8��t��I$W
��z�\����D�h&Ftl�a�2� �� C��yӾ��� |22dՁJ��$ත�n�K8����a~����nRw�������Q�������&���{E.��l���hZsd�s�@��b(�5���b�WbӮ9����f��a�HK��G!)�8���[�z|[���f��üB@�)���k����U��g֘]��;XZ����O��T북��*��*E�������`�Hc��q�9������#�]H����ȋ�GlyhR�jQ�_o�<^���|�������	:tҷ
����l��h��9N�.�N���`m`Q�K��?B��]9	�5�j�U`y�ɵ$S�`W��V�,w�ǟ��41�~E�L&��]eL>�:�F�]�B�����m�f{M�a�)}�M��� _���t��it_�W��F��5�W���̦�/P	I��2�ȫ��+����zrPURG�r4�Z�M9W[��"��u�Y�yo�EОW��&EAD;�����c�>���|gaA��^؁�!/M#������]�3��V͆1/�2ks�J���F㨰2��O�vQ���uF�O'#�x\ԏ���R�(�F�%��^�)��`�Y�=
��[$ª����S/"c!Ekա��,�Rw$�q-��\'�+��a��ثmje������QOYd��C�q���^����t7[5�G4�5����R��Hݡ���1I����d]�����{4�������/���O��xU)�+ i�U���� ���^n�gM�~�7W��0u���k�=nh�Ml�Z�$�jت��9���>�$ڑ.�ОyZ\��̀ϰI_!$�BV9��_�}�dS4O�;q���j6��E:a{��`��x1��E(�4ᠠկ��K���
!ݱ11�s̃[���?��f]㤤Rc�![i��Fu�_xS
L��h#�1�҃���u��&j��Z�ҿ�>خo]�ꛑ#DlGRi�~�#h"�N�n�["�u���L��a�c����nǄ��a�$�v�W��Ε^��vZ7���炶�PI2<c:>�y�,-�w��&'��T9�������G2�����TM�⧱YS'�B�qn��{;��;"������z��, �	!a�"7Jw}R(ns�rLˮ�š�9Y�=�%v�|���]bq�NUky�`d��3��ԧ�`g�� Pɍ�T�&?д��4�, �����m�YY��+d�E-FA�p>H����P%�e)<ܦ���	���ҕ�R"�����<6�����k9+���&D�p���΀��U�K���'�_�j1� 
����R���ggFDw����֙�8Q�c��ׄ�)ք��k�k� J+���3gjAA�!_��H���0۷_pu�!�� k�ʃ]p���pɣk M 8�w3qb�7�{[e-�Բ��z��u !}�Φ��=f�Q0��JM�JV8:���e�����Yc���$3��L�ۊwo�R��)!������o�w�
�+�����~E;xx�&�������=S��k1]WwRBi�E�Ӳ��^� �25��'��g��u W���?׺*$}���ԛX�¿<-u�..� ���N��A�n��E����2�K,�G#f��i�1����'9�κ'�[B�*�yݢj��˂%u���d.L�t�d@�"�q�ݜY7T�w�J@ԯ�Dw�9ʛy�Y�ѐ��V����ێ5/���>n�~"R��4}�U
�.�c��.�g�e�~N.nZ�M��k\��z��?%��#��K֔��#GXI�����Ù�	}�TӸ��_- �Mp��a���h���,��ܲ2�e�����[{2k���
+-��~� [7�ޘ�w��������Vk���ٕ;�~�K�SY��N\x��?˅�s�(RBo�#�ށZEq���Q%^	4��"���<C����]e��(�7�_�K.3�L�)�C36bsU��ܘ�fV��,�e�yuz?��
�L�o�L[�^�7�Q�<�5��P����&�2��w+ߢ�m(e��&u]��e�����osv�K�j���1����\峛�\.jmXPZ?q()��pk��ʄ�H�X����r�#Muwq���ң��y�I����I0�jT�`#c�~����Ϧ���&(c��K�Fq����Ɇ& <޵��r*���N4� ��W�����<�=�;*�J^��ğ���]�R�Dr�?�ӤQÎ�8n��1+:��4���W�31��0�*��.y���p%�?�%^�Kq�,�&
�I�����!P�L�7��z�I�Ć��c��T�t��8Ґ��?.Uv�Z o2<<������cc��j2���FՃ ��$�e_��lȧ�ökb7��:���AV������+�~�S�߅}�!�G������B {E��(E<��H�}r+7)����1�~�	�K�!HNx3���I��uHR6e�|:�ju.ov�!W�"&V5�:�!���1�*�ס��Y@"ڨ�\�F��1r����G�.c$�����J��Vha����{�4B�x���%	u�>&-�j��"�#EN�Z}�$ �W���3w�B]m����JպƩ�)����`�,�����;˹�8_�4��]+�1-ǹ��l����n�R�����
��J�Peӣ#.�
�%HW�IXK}S���KX7,��/��t���X�����Sp��=f����]l=K2Ͻ� ɷ�X!JU�I���7/g�	!m��+�)�j}S޿Dt��ۊP�9�vU�VbI�7��52CW*�� ��u��U3[ϗ�F�Z=�%�Tʇ�$[�"7�)"�ݰQf襸�>�4G��5m�}�ֵ��v/���)�h��1�/gX��y"e�9M�/L@V��WN�M����'x�7�����$�ʺ���@UR2@GMWA�$��6��p��i��6p���?�����AZ�LY�׽[_sڬW�������;�aŁ(����K�,>�� �9�����ˆ��Ѳ�?��o�J�)�Đˋ����o>��;_o��"��Z'�Ήr�2/]$D_W�Wmn.l����,2(�J2�l���&�.X�R_>G��HJ�.Ћ9Ε (__K7�'���p� DuF��Ac�='�MZDFg������΀@i����d�J�H�tF�uh�L9��8���	��)chmx��b�E�'����BG���1�.g��j�^^O';����_�v��r#��B4���eh�i����{��ӟO�N��w�8}����n3��/'6�oe[�OX��m�c�m4fI 	��Nk������Ȼ>�b��|�Q�t����
�A2��x4���,w����Y��1'&��{W��X/+^ {���C�i?b5\���tz>��e�wn�9t�f�J���^3S����a}�M�?�Ā�VZ� ��W��^�]��m��xVe>!b��>z��ٵy:K�BFO����;�C��`�֡���q8���
HKVP]j��3\�n�����$�g2Sg���$.��R�~$=�<�yD���g�Nm5ď��ͫ\>�R?4�IC�qq:����� �j��lO�S�BX��~de}ǪMmH�⻩!�ϒ�����S�ۮ�K{��^�h~t�/AE��!
�E�hگ�w�$���h7���#���G��á� ��}9��l��qg��*���{M�r�\�eS/���dK_��A0#;�,#��k�P���~����~^;��P���EtQ�,�|�Q R�DKbr��'��5�u^�1k�^�6kD�U�	2��ri���[1��y�+'F���L��Y;�BZ��ԌB�(����b��a��xG�bS�5������:��x��gZ+F�[�*ᴪ��ނ�E��x�\O�����Q)�=X����yP8��	SдS�����m��HK��d�YKNe#J�3�_��z�ݕ�bO���- Pw�~��@#�zdǬ!��������yO�����^bSp5h)��$�'��=	���'`o4I=m[��pk)��_:�;�v��F��Mu��K�N�3	0QXT�gß��wa���t��:N��%��9��g:�[Z.&�M���T]����Zq���D�6��X���Y��%B �$�_�q{$�	���v���ؐqȨ�<��^��z��ͼ�0���XIO���ÇIr;g��09Z��uI=��@���s��Pƽv�þtl#�.=Khf�t�bJNb�}ݧgp|䘣�QZf���.��t���ĵznVt�f �0#8Q!�|ɭ�B�0_�sE&��Mpׇ[��,��Ʉ�gS`�w��¼Oj�p�@�M�/�sz�g��Q��+��������{�(c�@��i�C�Z��aq՞�6O����\�q�.�|�<#��\,����yh;�R1�N��&:Fn���py�@8�v`(���s�������зX�N����_�&8Q���ϟ}$�~�a�*%h�0�#�;����u]=wK�L�/��yV����QP?h��/ڈg�f:fu߹��K��-�M��E����VB�F_9��Aj�4OgR�G�w�"E��[���Ji�@�G��
�M��P��9f���!~��o��ں�)�[����Z̾���,mRɤ=�� �.�ڂ�͠
q�!�`��C�$}� �����L�̹2y������)@<�oy��z��몠�+6k��yo��D;ަR孝�g�up؀+p�Q�$;��M���'oZ��*7#Q�Q��;9���k�U���I5�;���d-)��8�1��E�!,���&-�
��ug�K��ߟsV��'f�����a8�4�u�i��E�q5���p���\�ǈd���㻒��춳jY%|�Z��s���ws |
G���S����o�Y9��X'�������$�t�,?�(���hU"�5�Zp�����{_��ҐZ � ���i]vVIX���	�x�<�з���xj!nm03f15p^�L`��b�4->� gD����o��)���3�p@�� ���}«=�� h6��3_n��s�P��C 9����Ԗ}�&����ֿuI�������s�V�u�Xs�گ��	�%��{ Ҭ��\���l{��y�~V8dyk�^�@��B� �'�R���I�h�h#���gu�c�빟p KH�  �����+H�O�>`�論�m�e��2�{57;��iA�q9 �7��V��j��6<X����gL�!��}���|��R����wI��D����!�;A��j����l
�\���d���|����:�vx�@���X�T�����a����<�.N�W�e��,��P
/>�}�I8��N,���=�q��.�
�%�B_�����%v����M���M��� �M ����l� '��A��[1[����S�����V�T�䨀hķ�����D��)�F�,9+��&2��!�͏��̧�Ja���R�Ch���h����5�ȯ~T�	�� ��q&1�'WTz �M��Y��E�'!��\�j&n�Ґ-VXW,?Qf<4_���:���6��pc��c�u�|�	c�_��M��b���g	|u:�5̀f�Z.kd�=�-�۟�0�93$��������J�x��%��Qh��sS��'.�^�lJ�b�h�����s�qT�猩�9��:n2v��3(���<����7�}QW�-K��W�9	�¨{0���>���Cb�#�����F���R(�BN���e���ɛ��:�l�!*�6���*����_S��*o;�>w+S�VB�
c�I 4Z�`��?1Lr�q��d�;����A�[�#���ckY!M:"�tŀ~#7�B�!9:��D:H�Ԥ7֡~��TT�	%�����e�@�_ZE� LiE=�X(�zP�!���ʺ|�	f};�H�U����}k�/�GPLst�Ƣ"�ǽ�څj�7P.�3ı'O������U��y�9��`�d%P�!��x�x7�~��T�T�e-$�����pC[ֈ���w�����0��kb�L��O������VǗ�+=�����4))sKё[�C0�
��H&u	\Eւ�Bژ���S �FF����D�:J#�w��U>�sL�^*������W����Wt]`�_D����H��w����m�PLk��wtF�c��mv��껒F�ͼ�̪M�!��T��߫��2�,���RS�64�{���ݱO�Y�_�68<�;��R:����}�t��I���nn�n4��Ԡ�[��av�������㖦}�:������N:�:sK_�Lߌ3��H
��䃿Aڑ̏@7"���G�)�Ga��?��g�A�\�㬼��@u#<�~����C���콁�g���]�Br�8���m�T(O���}^��z'�0?���3O����v#��F�}���ׂ�5)e�-Fs%��Հ�|"��VPC�>G���������f��a0P�#�dU�8l��pSyf�]W`�mz�3Uۙ;�x���-Bp�H0�D�Gۤ2����|���x�Um�6yS?'��/;bd0~G��d���Tj�Pd�oQ��C�eRյXXm�*Lh��p�|7N^̎8cnM��$>UT�P�%�:�!#�e��3�qkQ���24�XMF��T%r?`}ސ��sV�G����b�T��X��4��S�u��b��^@n�h��`���a9T�)��y���ДFqm����GO�Ң̒H�B�
���V;B��aH����֋��dt}�#�f���c�|v��v%�J�G�c`v�1�5�Cl-�A�:�ϐ�1�c�$���&EF�4��:��j���1S!�������	b��(��Z�}Ϩ/��$��^m�O�U��	:Y;%l�v^eV��)���~�����?��`�us�?���N⹔X�쎋�h�M}�a���[w�t�.��7��#��_�`�%�7X�����h��9���j*�2 �Y���ޛk�,uN�#�>e�Q�(p�5d�B��.E�	��&�l�>o�2^�On9A�?`�r��w^��8]��.S�tɑg�f��.�U���Q'��ݤ�GZ�+�:�)nG��-ʣݡ��(�ہ�=�M�]�r-:=�N�� �h=5���d"�b+���iP@�	Ga�2߽�y!Ԏu4ش����Z㽹$�є��)��
�����+�l�:C��?k5β��uo�:��.��I7d�����Ӯ�1����'$m��#3Z!\���{a??i�y抧I��,߭R��6g�[�wǬ�62A�Ĭ�O%�EZ]�i���a+���M(��=g�ܪ�V�]K���T�n���;�߰��� Ez��J�'Ӧ2J�1������r[����#�"jA��p��l|@��Y5ܐ;
~��,�O4H6F�3��3Û�+��J����]����9Gk��������ZP6O��lZ!�0'��Ӆ<�uԎt!p���9�N�8O�p�����T�nD#{Ҏ�� a5e��e����-O`����������C�mY�i��BG-��P`�m�>�b�#�܄Mţq��M��R��3E]��1�l-V��'�vi�}8MA�7J`.ck;��Y�ZҲ�z��©��=#[��W�Ey�5t���ݓɪdF;nD@��H�@�Y\��I��W�+�ȣ8a�>�Ǔ����@���P��p"d/_]w�����}Mt��3ׇNI�[�Y�o�'1
�٬�i	t�${SK�^4���e��B��g�+�g��f�އD��j𬶪}*���_W��xSV�UC�[����y.�;ˣh�Pb�=$^&h���w4k5(�Z[Y��7ɿ�K^y��~��R���ZK2�x?،���
��!(�5�#�R��)ʪ�J�sG��P��{4��Xڎ=�Θ����ܩ����,$�(�Pw?�{������Jih%d:iE�K�o�z�ɷ��^D�;�;08a����.�lk&��/�]s����Bױ<�7yhp;����(�[y�������Ek�Q[��'�>�dʇ%,�K�9�#Y>[��򯇀�v�yЬ�i>L��^�~�����ͼ4>o�&�Nd�Q�zb�Z&�.Qz ��Z֪�:���K�0Rs�ƹ�LrC�9Vm�;Q�e&S�1d����������+@�YI�?t�xˤZɂ7���%SV�(�pw��N���v�⤾��C|���F��^�cLk6�����mG->a8��}�;��)6/��Ct�*�;��0_�f�H��?��r���Y�μ���#��癡�=P.G����YiU7Ma�xO�YxK��%�v��6�ѷ�J�0���{zl[tdo�q��C���u���ֲ+jD��o:*�E�ܥ .cW%�����M�m���\���� ����VM�m��x�+�fS�w�P�cO���A��Z��cmykq���9��~�/X�.æv!�4y��N��:��b��Q�z6�Lq�<z`��'	�mɣ�DA�5�Q�bi��p�޾���*��E�)�0E�����`c�9E�U?��xG�Y1~Z�[�Ŗ�RD��H��d�]����b����}H�I�@܉�p#�X�Z$K�P���0�N���"D��[�P=1_�Ӳ�%"]�OQp�%w*E*%OZ��Y������<��n bsؗ%���S2���&��zx ��K-�wp�B����5��d:�c�j����b潆��]����eF�Ba@����#B-���2?T�f�:_M;��f�>'FtB�� �k.�m��H��V�+�jmI�	�8��2X]�
��+b��T��K^XE�L2�*�j�H�>����D&~�b�]I��9XߗW$��H׾kYa�B�4*��7�P�⽂I}~e2��U2p��7�FBa6Y:�u7�7���)(mR���2�>5��7��\xBa.���+�+��m�Wl��h�v�9��vsշ��'��[��b�,��&^��TF�3��ޚWַ}jI����Ε�g ����W���،覾�a�O�O��XO�vC� m�dD�0g��£�\&;����
+^b."�O>v�@(�)��@�/^���2&�ZX��Ϧ�P�7��-��`Xq��75����o�*��'�[Rl n��	؝LD�C��7�"TJC���8�ӭ�Y:S��Z��̒	����T�ޏ�J��8h�_�� ������.��e�j�g$���U�?� �X�:����4�J����O��>��Me�wA?T��U�~��Pz�UG�h��P���g��UO��Pt��)h�,[�9y���a�@F�� �yY�(��t�ȟ�u�<?��1�U�T��;ޓ
Ǯg
�]����C�7��6���:��q}��.�A�1L���sQ��7�`��93go��⪠H�"n.��4�C���\X���\�����s&�mi@�k�Gv-Y�
�XD��=�e{���4�������9�T�LTkI;�<�o����0m�a����B�l}q��G���u��i�'� �J�O���9��B��"8v|<��tLE�,Y%�<;<�ӛl5�_r��j������|}S0Ώ���G�%�VY���8��Q�)hkr�y�P��r:=�+3Z���CA� ڻ�Z�X�e*	|�ty�5O�g[E줈��Pmnuif��V�J�D}�՞n�%�_��w�p��n�\`i��>H�%�H���O��(]lxU�MN�����T^�SL�a���ۓ�x0�P��
�� ��!� 0��>���6��]��Z�O�s�����3��׏2����&����E�H�N(v��e����u��5
��;��Z��V������f>H	��`����_jjЪ�M$rQ����o	E{"�H��ʜ�o��ses�o��4���bX�[��kT��nC�q�CŒ�>r�_?/��Y�r�/k9�����WY޹F����D�\���
��	#�
(�$�0�+;����W��h��{	鼇)��&ah!"������l��@*k��T��2?0�;�$��!ӏ����(�L����˸�۬����!�kDjH�R�'	OT�k�'W��e��F�n�ذ1d,$�����,B�;z1��n�4�W��/J|�O>��Y�2tސ]l�����&���ߠ��s���O%0�ϓ�P����Q��Ë��S������|KBu��w����{8u�:�r	�y�Sʧ��5���-���dn�/bV'ٌ���!2_��N����vK�[�t�чD�"s�K�C�@��=�,I=\*�,����F1[��1݇�(�4j�f؈��:?;h��d���Č��\�!F�H�t��V�@�m�S�}���Lc6)��Vj���vXx�^@�c�-k�i<Ǜ���P���g�K�p=tz-Ⱥ����>{��Z�LOa�}����C��L��Ul���̑X͏���#�!vU����G��C`r�e��P�ϗH��Rk b�TV��@F�y�[�u�Eu���~5-�h��%T�F��|��"j�l�r�"�e�u�Í��?�(6�8WO��J�@Ea�8f�J,��tb�/��zrO=�9�x�(�����8�9�j���,
�R�ځ�>�|J�^����WLJ�bm=���-T7�N���9�@�ެ�D|�䄂g��AD����0�7��㟈��@��fEѴvE/��Q�b�I/R��u�jq�7ˆ=�mG�	��A�
��1"b�X%�~W�Y9% ��;4�W�
;cĂ�\�<x�$�XM��n�U�P,I�ǡ��5۫�o��S�q����/^�	oCuϞkU��;�
�$�����w 2�-����͙������j"c��T%�v	k���#�\ׁ*-"�
kZ>r�L��t���_��s���#�!dt#*�.�\+*��؁32.z�R�p̉1��M������`��{Vl�$��G���vʘC�?1���C�7ېv"�f����O�[��X�Ǻ_t��D�Q<#pb11҂H<�>���ş��ۻ�b��	�6�t�,�0~՚B�2��pM<�4)Lϰ������+�!��쑌 ���4G?��¾�$�p(�չ���5�MT�(��P�h\�;�S��TxxW�Pz"p�LF�|��XX�3���4`֒�:B���sŘ���4�-�(D��R�S��E�Z.�iot�`"�Ƣϝ��R��{Q�e� ��id�)� ���¢k�&�3s�G�w����mN�A$����bi�1m1�
�b;��s��%��L^��틔��,�o� �gM��&�.���B�[�ħ
L�)��1�(�����mDl�k/X|�+S�������@UV���n�T,Z4�b��J�����FE/!b����&@9�~���nD����r���@��I�:��	$V5�:�:{��l]{m@l� �|��px��86"~�le�o&�g��Q�����@*03+�S8��7�
[}��:����둹QMu]/ ����P%(��|N�f��ϯㆪ�F�O�Lf>�\c�.:�+�;x̀F}x�|�`!�nυ��8��7i|~�K�5 �?QzνN�������#R�R��~9콆�O��_QE����a�M��<����bz�[��#n�wT��(�[UK��s����6ǎ�'�l�e�{^C��2�̔������LР��V!�}���
h�>0+� "ɥd���9� n�'ɺ*ւ��C�l��҅�%|z̀af�ut�M8ݹ�_7�IQ�	-��R��D��r�U Y������v�Ǩ� O[�Jcܹ*|�E����u��rHK�H>�F� }�)���va�YBF��Ju�7�:1*�s�,�:�V���etCO�i������.^]���Pd�K��P)�xN��W4v��;�m֞���'c�;8�nP:0�B�ڷ��v��G�A#$��L�"�c���1!��)��5��z��0a��Ui�������ى�5 �H=*��*�켔�C!�1���0Qls-/��n���[l��K�^�۠'|��S����u���C�G~��������c�y����j(n�>���g*�� -�� H�"�u�D�{�>�!�A�W(����;ܻ��	N����vLW��¥�h��j�d������62��g�2���< �:p��A�W�?��%����c������Ռg�#pw>��j*}�1*�!�%{R|{�'��(�c�����l����@��7�[�Jhi��wgr���]�'B�=��4=�|��� �w�߄5���/`F��=�a� �53 {QTر��`t Av��po�E���W���@�L��Z-��4��+F2'Ⱦ�*<!�/��I�f��dK���D5�5���R��,�N@��qOb-�e�?�$ ��u���0�!ǐ��q�,�+Y3�� �R}ۙ�c�$ًۉ3���o|���)&�ӧ��C��kL��E������V)�͌W3(-`�̆�g�J�֗�)�x�3D-ȿ+�)[��O��/��j��,���$�es?s��)������������!iyx��:�'?���d����[�.�
����d�]�U��Љdh�U RPO��׮�=Ew�'�E�jLrPO�Em�9���[�' �ZޛP�q���U����z������$�4\zC��9��|."�22��Fe���������f�[�'x�K�c���G��������e�5��Nz����b��f�V��^_ݐ�P�9��������H���lc�I+_j��N?|\LݘU5�)�S>a3)@9T6����a$@���,a9a�"c�$#6�O*5�'���n8AiIn|Ȏ�YM�[�p�[��4�nVI�31�Ҽ�Q��h���^��2��+��'$e��R�eL��d�x�r�����k�}E/�>g��\.�5�&���3_gy�Ă�!�� =����&W����Q3F�-
�x��I���)��og�B�T�S����V���bi�2۝�gz��S���`fl�0�a����	��TVY2�z��!��T�1s>(|1�~����:@Bx��J*�+y//U�� ����9-G��(s<�/aF��Mk�@x]`$A��`L��'$\
���ӷ(��:x��dl���%n� =�p5�W^9t1�%Ub�T��S�~x�3�!���O�H�:f)^����l�.�FŢP�H��&�bP�s��{A����ZTN�� +�P9dM��[��Ñ��!��Ɖu3p��Ջ�F8���|�	^J1�_}�S���G��gz��w#�K���|#�$h>j/ɜ�(�ʵ "�@��:Z��-�g۽,�ƌ�_��b⢘��f"-�f[ϋK!������[����iH%K(m�Gf�]��^�����݈1�u_hn������RjO�����IM֮�or����vh���
9�1�+=y��o��[?�ܝ��_i5f���j�ZG��I����Y��S��y�g��4���+
�f�NH�l#���/?�-�GB� [n�C�������z��p����E|C}}Ήu��}t`v��$�'��=e�*��\��(pEhZ���R�(w���O��kT&�h+I&������7҇�/�˥�/6#`���
��w��?�7�̓�Ȏ�)��GAD��\d�rǍ�)�('-ڛ�r���I�G��S�	�6_S��� M�3R̗���%��1�L^�ϳ�:�����Shi�	M��fG��Ix.et2Xujb�Tle_���C��`2]�9��;�u��Cu�I���2�I�h�y��0q|���%�z��OŨ�A��瀛������@.d!��M~ ܛ�>üV3gO�8�����S;��G9n��#6[%9�D_*X�Fw��ӳ�L�L�iO�?_!��Nґ��r:#��q=ln$����~� �v��5�n��S�$&Cy�C��7����2n�ZǓ�M[��آy�k������mw0���w-گ�!��vGͳA;��?�*�	�hC{e�������B��x�����Q����2y)�,�`F�i?W�6!���?�*4b���B'@�]>�e`��G.ßv&��]d�Cx�O� M9b���C�N�Bc�n*0�"���f�L�|r�ɥA�MS�L&L��h$�Qs}�[�ܧ������7������(Q���8��~&"�a�ƸTVH���}��V�'-���0�L�+ Lⵡ�ѓ�	2k�̄�4��� "��c��g��2[:34@�M��<;�o�,2y`�mf6�Y��4�{�(֧�|�����7�qelw�A��X=�_�P
q"���H���e�^A�/�EV���q
�^�@��7�Q��AI��)��N�8{�r9,jwi���N�P%��ɹF�4�����U�G���̓���4��'��/��r,/88GUk�`1�]��V�p�@=A>ajSg،i�����-Թ%��kR��aE͸�����N����b�4g�;e.Gޢd~Ht���m����?쪥�>���v�,���!��EU�3��:������ʑ��k��b�\�=3�Ƽ�AfAc" *�����Ty�񟏔ɍ�*$1>]��jj3�����$��,�t<�B��P�eq���{�q��Q�rg3ãq��B�螭��؊'��
F���b���a��Ude�Y�Q2�����kbϕufiG�v�+6T{=�QJ$ǈ�}��M�?6"��LL�A�ܦ��oꝓ�]q�-3�7	&/\�F?~�	~6e�(P*%%c��2�iQ�k��p�)�[��F[�Jx�}�v�Z�
�ԋ��}��lҔg>���b�2nT>bZi���H{r���Px��YW�u��5������Ģ7�H&���	g�.��n#�^������Y�7���C��29��y��'⩕�Fb��≴��a��isϬ����y�;��7���3sO��ߵcP�q�cyl��i�%�"�m��мp��%��!�ez��2H����I(R	#��6H�Ƭ	��w�o𣞵��U=�St�"P��O�vcZ�X�R�H���K_�
����Y��u%0�8�߹+���2K�/c�q��Qu)��k�Z�5��k�
�梸%WJ��P�N]�@�rD/Z��}���i��b�4d�[�X�fg,�Z~.B����g �:d�`��-���U)U(��-���!I,y��-��i�G? �P�Y��X���MIc:{��*�˗\�*�����j���C�xJ[#��V�OvY_T4ׄ�h�סI��~l���}Y���Ս�:J?���`��*�c�+����Z��b	g��A{/����#_��p�UZ\dh�@k��w���á�féIWvNw�2�&\�$� ⢻�L�{����/?o72MO�})og���r�Zf��P=��O��f�#Iͩ�:����5���8�^��0����_�U�{�t�UH��$����G?�E98-H�P��(�ŝ����DK%�};Cnh�^C+
!W���{J�v���7,@�"&�"�'�H�JV���F5C�]��P��^�`]�"����ppܧ�:g�M��/� �U �1���D�9��^�6������I �?+���o�+�v��W���h�QR<K&o�Z�Nt%���%i+��lj��yo.������P�o>&�"(��<kC���O�5P4L3���9[e��D�����fS��sH�M+yS,��U��T��i��V�"����V�����?d%��_c��W��uL��Lj?�7��9�=}�D,�j��ޣֻ��"P3�Y8E�
)UB�����M)���=h��<k�_�- 
}lʕ��Zt?	(`H�Z��D�"���4d�܋!��� ��M^��Fs���ln���A���*r��;�\S�bGܥt>f�n�k6Ʃ���Qm��C�ǐ�j�����]�99���)�"�����tN����=���s"X(u�3��*ۡ�x�������N9��)*,�]�U�����/�}�O�ɱH�����k�%%�K㪞.y����!|�CBZ�Q	�6l'������ Ҍm&���� �3��Z���MB��=Ŵldsi���|��캑��9���0�d��A��u�|a�۝p;H��� �^Om٭7ͮ���H�����<(�"�4A�1)�D�a��L�3��Y�&4-<�޸��l��t�����QE'��B�������H�D#/
�[S��E�t<���Ÿ́�2���y�w��p�CcN��u�΢�����ڋ̖n�	YK��9Z@N,(�L�(i~���Q1#�i�0h�t�}�;,�؈٤=�E<�y(�Y���F�JP�6�Ԡ$����#=IX�Ta�6�\��J�he$�e|�=Xw��]��-Kߎ���~�*)�w����/V�\.1
c��X�Q��[9��=��":Jo�</��:��{H#��֯����M�xg�a�(H�yTak��]ݫ�Yz��.��Y0E����Û�?nmЍ�w���+l;�Z�D��O�:�Z�"�l���K����#�g9Ѽ<��j�+C����CU�#��3j&K3��9�Sx��Z'.l];?�#l���J;�P��3S��eѤ�!=hlB�pCʌĜ��m��-A���ʒq����w*zIq�@f2i�R��I(N�)LF\h�v���o���AԠ�qL�H�ǝ���J��y�|N�ʍ,�����=�j�4�u���(�����	�N�d�����RG��?�����f�4θ��-◇�{X�����R��5K�4�.g��+Y,Y�R��g�����s���߾�4}K8��v�䡯��*H�e����ʬj�Vk��/Z׸�{|���\��J���@)Xm/������;.w�9����h\ WC%�R��1�eSԛ����H�Yx'O�V�	�D�ږQ��%d<�)���]�h����чƬB�[M�`��*��Q�w�1aP��Pf�ˤ��L��L�$`��)�.P�B�g۵��Ivߞl�nft��Hp���E�ښ�rar���g,������6l>���pK�2�,���#�x�O��%��;]��֯��6\$���Ң{E;+*�v�K~�hn��(��)���������Z)Y���l06u���;���,��Z�@���[���h?�/<f�K".�âh}������>�R��
W�F�_5T��<�o�P1YNTs�@�� �bf71��$�d� ����7�=* "D���*t��������X,ry9�Ik� �;h�$��W��2�y���Y�%��_7���h\��X��ۀ^�G܎`~�g-�6�$����S'$Г'x$�
�{��G�*�~
���B��@�\�����+X�J���T\` �on#�ܺ�J�Xk~������ǩ��_�7�oM�v��"`@�_�*�'-ԡ�,7dxs;OT��.�0��<��wB p��S�*����,cT��\��*����T�eea1rj�,�0c��Y�g>|��Ã�RC}��ܤ��P����CӍ�޲�Kζ*(��-�ukԂ�e\鿞�D��+/��g���c��a��{.��du�-,�X)U�}�ie`�=c0�蠫h�^�)�89�*��W0���������v�[�(���o����2NYF;�p:�y�(�􁫓p��v~@��X��i����������&qr�%��Oת�5n\�W�}�	T��y��In��.`�U�*�]5͢����p�0yd�X���P��6&@�ĺĒ9_���Zc����x�r�	$W�o�!���q��w,�3b����dk���g�`Y�SP�<�%˩�IG3�S�=��;IY�T�����Ľ�7�zP�jQ�;�H�*6�y���r�!��ะb$�R��ģ�D�/��{����+���h���	�mvQrH�?��H�,k ���T���5�K�������wu�@R�S� �E�Z�×����oX��@��c�*2�2>�Bjc���Lc�%�Eyg;�Lm�#h��|R�T �1����o2�q��j�\�'��h���ΩԄ��ޕ��:[9|��;]%o�p�3�:�Î�j�dI�����o�rB�p����lC�_X	�ԜŬ��e�V��o�u��K�yM"�G���·���P]f�r�~��e˨U�;q1�/9�p�(	<W��kÆ�f"$𥞃D��r���[��o{�Cn���(cj�I"^x�*��kqz�
��vv�.Q�-�da��Hk'h�mr�V2 @�3H!��iO�5;��ؔ���E��M���o�i��ơA#�P��J�2��I�id�E��cG��ovHI4X�(�����z�=�ǃn�$��.]+����}�U{���pC���^��kߤ�k��Ԉ��EaTALI=�V&�] %�;L$&-���6j�t#X�Zr��%��NQ���ȍ��1�������B���6F�1c�\����Z~gT}�dc�|a���M��%�K������)��h�L{�SXfCP�$�ۋw@w�Ð�U�ÿ6r�Xu&t�XM��v�{����u�}d5�.|4�&���Ƿ�{��ǜ>�e��R���j}O�;��vCr�]�R^m6��c�Ã����g<�]��`ړ5��	H�I����l' ��7	G+I��Ꮺ(�9v	�)XRwUk�_DȰc�����ovF����rFc�K*��y�/�_,H���B���a��� 8� ���~
�!x�,�<�� ���(����M%H_r��g�&����'�̃�)J���`KM]��^VĬf�Vfj(n�Cfr`�w�˄75��A��c7˷�T��R�6O�k5�z^�& ��]X�q��f���o�� k��Y��g�����}�Y�.��9�śf����q�f���3��[,��zf�M|6���v�?���5p)�|l���� �]Qi������%�H;M�i7-�vU��ٰ2�9�J�����M�O$��q!���M]_�n�f��m�u"�Q���{<4�XniwV����<�W�1��!�����	������oH�N�i�[��?Zk<H�G]|Z��y�f���A�������M���E<}9C��Q;@(�ɖȈ慘] ¶%}E%=�����2���nM�#�+�Ɍ�\��w��q��.�Ƕ���4�ʙ����%�*�����|п�)f@�4�ǫB�+���UMiL�׃�v�s�g�q��<:����8��Z�4�غ��0	��L���k.�wQ���0��IVTPn�z�{��<����	;P�d���Jf�v�(�t�|~���i���it;��mQhP�Y���6�B�3�s����4(���{f#kA�~ʫ.����̫�Ż�dkk:� �q��(��[�οI����+7�q��|��B?��^������$p2�N��ޛ���Bk���
���y��?����SB#��۔0	����p4���Lr��\�JˇI)�2�o~�x�IX�LFW�R�o���j6�>�h�R��9r���\]IK�w`���ǎj���t�Ql�rfwa.mFz�n^��dq���zn@Z�d�W���@���3ƫӵK�iCܛ7�T=��[��.��o�Ы(C\7t����Ӭ��&���f�2EdKv�ӂ����y�M'�ΡT�hBtcF�]q������E!�{#_e�'̼wi��U8c���x�C�,����'� �5�r���њ�m�2��x���/��\6E��W_U4�Q�{���>*�������+��,F ��%���!��f^����t�?qk��'W�o �.U	E��Kp�Y	X���n�Gjc+��֯!j��6��E��W��ڠ�7�����Qz��'q����1���7�_&�b���}@�q˫�о�>/���,��99���|�U����u+Tx5��[2v��V53�/n�O2�*��a⋼�n�DG_�������y�����;hG��E��%H@q��2���ƔQ8b�pn��C~��b�ȗaW�C�o?�����ʈ��Q(�VF�O�h��/#3�6Vw ��N�h����*�'t������O,!婫ۙ7��Q��O�`��k߇c?tHP����U�T�!���N��cؙ�β���,d������~!,�H��ݩ 0���!9�������xې"u]F��]�拤+max��S�!�">\#L�?y�.t��V%�������fM�o�y�^��d�fF0Q3�D�\iIC��A�	���{`��OT����H]�:�����՟Y����ő�23�f��_�M f��ڊ�������?�w�0
��H�Q�Ôg ��r�K��Q����;�Ϛ�v��T����j>�"�b�	 �S�f\i><'L,�OӼ$�t.5��	�����MVM��\�0��k��1���_�&�!ш�����e*���l��P!�*�-�FB��Kt="U�R�k%�Sz��ݨw��<�u�h(>��U���F#X_���A�b��s���u"��7z�,؆Zx�BqcEq�����s���xw�?]	UH3�}�^v�+��Ȁ!����`B�W���ygr�"�V�4�h��b`g;TTB��{���ݲ\���3����U�t��L��gOW O�i�zى��Ϋm	uw���O,�l����ֳ8���܄]#hA6~�~,����]��$ 8'1~n�w@j>�E=�}��0
F���Yu�n�p�R|���@z�'�'��%S���aN�K�{����N����{̈́ �͆
�s�{��g�jD�lE�*�:)
A�V��t����(F��
�ҪB)a�����
�:4��z���DΓ��glN��}�>�Koo��EwG2Ɍ&��S��MT|�NΔ�`-e�{��	���)�2}_ ���(��͹��|H=Ȟ�bR�DP��҈fN�*+;�3��V&9|��T[�@5����ܼ{drb�n�6��4|`����c�-x��g-�!b׽Ĭ6�S]��� .��<�6�R�E���<[@AXD&��Z���tV$��8P���&ZV�;�k�ׯ����I�^k�H� "u�����2���4�[��J��?�/��IKB)Q"�Xc]���1�"_���p�o`��R�e�}��^���A��r��b��N~_b�40�<�Ϥ�ڢ�߇w���Q��S���y/��\�"/���'�j�,
ܷ�3$�梸�!���Մ�]
rR���VY�9������y�>ua(T�0Z�%E�x߰�?��鏇�A8�G�ب�^��-�;=����i��������)�P��]{�_�t�����\�GTj�c쟬��R�u���I����B��Ʉ�q�$�r1驂Q�яw����s�������\�l��������\j0(fF�j�j*o�Ҟ��EUC��a9��S0�éx����H�*�#���Ｙ#��Z=�t���ڜ}�2q��h��s�{��ɭ~F�������X�y]���l
���Z�7�j�.�Y�E#�@z>R����&pkq=Dd��GS��x�W�֝��wĀb`�7���C��)�Iˡ��-�0��D?@Q�Qk��Q���ٽ����F�A�ۦ��Dч���D�M�ِ�E�5��d`��Paz����3M��P*�7,�[�0��۩4�e�χk��G!}�×�1
��Y�q}X.EY^��N����o�G)��>Y�O�l!�{�r��I$�YN�),�p[� �v������e��s����#��yI��P=Ms�򥠳��R8 s�/ͻ<��7:r�ժ1#xJ��09�s���tB����)�zn�Hk�&7lʂ|�e<�bZ�����r���.� ��V�"b���� $����Dr�t�u�����h�}�h#�&���tI���3��G�{�2 tf3UH��gf�L'���x"~�I���Z�,~xsg�֤�%E��>o��ܽ����C�/�����D�Zx��u����J�9���do��m�v{~
��S�L�h��O�Ƅw�x�p�N���#4�r
�M���I�s��.;/c�[=�xR���