��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��s������\�Ἡl-�y�f�����f� �ѕ:�nA�kb-q��_���ѹ(4�dê*���7��N2�ɐ��+ٞ�4Y6Mx�ejǴ�y9�����=���D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6��\\�l�����r9s��@'�k~�{�<���y�#���i6`#Ɉh:^[����*`��Z��|���z���N?`q_���ר�Z���FLe���Et *�mk��:�2�|��S��1�L{��:�;��?)��/os����$I�G��S�Y�a�.ڌ �|\�E�7��RH�����w[��`�d@�<�S�쇦��y~����췔ڤ�8��p�%M� �;�.?���EJߒ=6���o7jr����SG�C��,��)������ݍ,�aj�� m?N�L趎�i�eb�>��Æ��򲃁Z�7�	E�͓��rH�s�&��7��_��
e�F��H���)�W�g�l���[��燸TɆҭ�V�{�Σ��G�kx(�}L}j��"���*���A������s!ɑt�`z��t�ۣ@��� �f�wA�4��A2��rx�Y���C+���:Ѿ	w��i���5p�-�� ��Q�tMd�ei�oX:���}�\�C �\o�r��Dr�����dF��]�(�S��ş��#���ᤝW>Uu.σ7f� X��d�� ��OL��_KT�2�&ӥD��OY��f\K>�`q���r} ,���)(���q.}�3I��'38�X@�S��lN���x�Ԇ���䩪��J�sV)H���1DJٛ����+c8�{R!�M�4U�2�ؒ���Fg��U��,ޔ	��A���ޤ���&��� b�,*�%/���@a~hw��b(���'6���� ���P�1D��J�t�K�]%���l�4�ڹ����c})�wk ^�|\eѰ >���Sg9+R�䫍�0�̐�l��˘A�u6�N���,��aMŹJ�$�����H�>�:�RU��*i������ ����H�&������{�%�3�/�X��\�T^������y�YV/�!C���l�9��GSz a���y~��'>�ߑ�3E���ȍ�5:2�Μ�C@�Ǫhۊ�z@ˑ�A�ϲlk_�=��"�FA���P!�6QLN]ΆȴE��9吉9�������q�%��|��h?sI=/-��b�gh���Z���7�P������,�n>2�mƓ3�=n�}&�xAkT���γ u*_�L�M��cl�^�,�U.57s�B'7�W����^G�$���>���#Rk�Qy��0Q���G�|�O)d̆F�T���Iw&���ޒ��A6���9�C��<�FՏ?�Q-�p�#O��в�Y汊5�v��&&&�z�
1m�Dܭ/B�P+[�i�t8��<P��RЍ�)�5�������ȔǷ%��-ڱu�jQ������wN��XU���Tϋc�-a�PS֑�~i��i�\=�j����˂f5�<�3<-=[�7��A�ݯ�H�����2=���"Pl^rw�rU����b~�լ�b�IhdS|xa��yn�#!���p���_b�Gp/<y[�a���BċU٩|��v<�9{��F��g�җ������.5F����un5�����|�{���� W����⳻*j炖`j�ϲ`���\����vբgo<���{c(��TI�^��Ҟ���6�1n
���h����§7D�(�G�flx���ٲ�;J�����CKaW�g+5�������Yƚ�����(`(_j!Y::'�q�?�j�G���27�.4�O}�j��y�"4�/0_c��õ��0}�4NƜu���S���xj!_�f0��ʥ�3R>�y!����5w�u2�������7X�~�ȧ��+�q�3bQ�)�\�v;�4�qm;��|�lgײ�)�v�G Z��iL�[�2@Ԩ8�W��G��R���Gy���I�[0z 6h�ms�Lu����R*n��tH��~��(�3��?���Il��w �.�wrV��&�1x��|e���e{w�:)�(d�;�����^!��*���\�7����� ����)ݧ�z���&�����d뾒�1"c�ssX���f�G���	�����^�`�T�PEi�W��5�>�__�`Z��I�8�E�I��e�;��\��4&V���-1�u2�T�'��M��D �[
B�2L�&�8���C�-����$�qD��� v~WFi:��c��{��	��.��5��AP�����z&�R��כmz��u�U}9�쵳��0�E,Ol����Ṙ��{D�=����-j��@��@�2@�hs�+�1���7�Gf�9�<�N��c#.�,{a�G�҉B=4�j�^u;�c�ȹo�I��d�>W�XI��d��K�H��K��Jo�}�=�C��>`��	1ߦr÷WgosyW����h7Fn�}��^�"�ax�{�w�"$`�E����g�uz�O��/!���	գQ[V��PI^f-�FZ��%N��%��>4�OrC%:Q\	E�#��v���u-�UC�t�K�W� ��s1p����X�*�i��Q����K��8�P.)[W�"��-%p�s|�\��Q:�����A�1�~p�D;�������zDz���>\���ĳ
����Y�D'':��'/G�u����$���@4X���	8�b�Ȇ��U��s�X3��Z�0U'�fZR	�y{x���e�����l����u��fA�����c�Wٞ�|��qx7GF,Y�E�\7?��qL����~���D��ۉ����}�K �7"�Y�ǟ@I��:[Bϙ[��S��Kn�����)���l@T�y�nͱ��|��p���U���p�1E$�F�N@V��.E>{{���Ak `��?נ���~tj�2��(���s&JFp��<R5����R����Wz�m�a�'�{�PקD	�$<G��3s�0�n�=�"�`���sV���s6c@��f��iJ�����������9��ٕ,s�ZO0ы��w��_)�Ǳ~E?����m��J(,�q�F՞�L1	���q�r.�h�B+�\4�l7�l���p"I8�5��1���9W܁6�Ş���@ȍ�F�ʌٸHI4
m���G�$럾����z��-�[	h����K[�E���-o�_<$�؀���O]I}YuB�743he<��!�q�w���Ӥ���Ĩ���E���=��i��N%��el;�!����F@8%����:�W���`X�����=����̀;=eNB"���];憊q'oXj=ÂhK�����DV�7 �u*���&���EbB�%6��i���i,-�U�Q��뮭b>��ؾW�u���1]�N$���÷nR��U(�S��?|ӎz}�P��*��,T�Ĕ,���-��t�5�
���y2;��}���f����9��n]�)tR4|��TB9@q�*��Cx��R��a[��ٰ�R���:D ��:dIv��ivӝ�<�����񂿀^H���ac1�C*��
^����3�4]�So���!��Wp���0�h3x��v�ю��T��mĊ����)����(������O#{iG���@V`_"����>��{i�����I,OI}$�_�>����^�.��oKU��`�09�w�Ea
�Ƚ���|1��z��P��OL���ʕ+'�
z��6�bc�%0��9CѬ�\)2�}�Yh���3r�c�<�ʝ�J֑��6x.Jg�*�+�c[�\����t�|�<�I���\M�*��Q�0�8Z����7T��j�Ӯq����5�a�e�cK�������4����oS|`��z�<�ډG{�|/e)�w3�ͱ����
�udu+�YN(�.���~�%C�|�<�pZ?����qs�`��*É�K,�j��sV<�ɑ|-��@�(V[R�6�-���;7�$��77���Z���8��
��3$ݽ����<�����68.q���q�i��BG�3�9Di;�[�����c�7�*)�-�^��V	bP��e�i�h�v�w�UY���s&�ֳ�l�a�I��,���)����f��_Oz�!׽pG�����e	oC2��~Q��0|2���4T���{ C�
Yܜ��l���Y���L!�[��&bk�5���(,6�"����	�w*6��q,S�D-pu ��Q�<T�װ��f�Q�hI9<��s�.��:&�Yk�i�d�t��kC�PoJ�\n��-lɮf����^_MC݋'��`�{�p��]W�)�\p��\��و�EA�8=�gƤ���*2��)X�$��*i�y0hp�ߪLK=���6c]��Hw�E�H�R�3DWCZ3h7*"d�I�E��lX���"�p�J�O��>����x�8��Y�-|1O��5��� ��?O�:����6ˮ�t����G�B�X MG�-�#�.��`��~��Q-�k�����R��]$���^W戮�5_�S+H��SK�����#µer���u��FZ����0a�bg��՘��1&%h��tz���&��&8+����ˈuC�}��Hb_]���j�S\.�B�6�P��G�s��ٶ�L���l��5
����4�t���W��B�U����Kpg�b��8F��ҊK���5ݔ>�et�P`��,�7�ɤ�i7?ǂ�D�²P; ��V�ցV�I��%`��D�F�zp��		���
�}@��\0�|���,sM�%Ox�[;��?b[h�v�{y�L�s��E�A�-��)�^�V����﵋�/���P@Z�0e�z�9n^h�O<ц�6�x�-�VDlhe}��i'>���4��f�A�U0B_�u��9Zv�Ϯ}�%O�����a��kC#�馌����E��Fh�A{��� n?������=K�6,��KM'n��J5=ѯq�G���u����H��� �6��Ʊ����|l\×{/�[�������ʐ9��o,0�f�[�'t�x��3^f��#11� bw,�U��Aq��\�qVC��7�(�dy�pZ(����Dw�j*����=� ���,xpm��e3�̨��^8����G(u[�T�:��D��:S��]��m$I� :l���N����SE�$bW��K��c��ۂ�q���p�@wbK]ș���q�"�D�T\�d���w�����H
Al��n� ��5R�a,�J��~�3�8�'�ɋ������o�E�@K'���������@�t����@��B޽D�P�Hn��2�KH�)���v������E��5�&^�^�W?�B�'�xp�=���V)�>t�h�f�n��Lf�� �Ŀ�~�k�V4��"��;��8܈1����n8�ˀ��+�wX�掭�]��'�We��'&�%z[�uq�j��ؖ.�����W�>*�c�mV�e��S����dկ]I{J�^?L\a�ľDty����K�?�}�o��"&9ْ.L~��Q�4>�K��KU��:&� _`�h�F���T���ܗ)�B�V��C !S�ָ�N��a���?�����鰘�q[s��4ր�f`��9O-]�6�{������D���,#����}��ɶ�dchgB��#���
:(aeZ~M,����r��G.&���La�)���%��n^�N�Yw
!ފ?k��D�R�L��ޜ�ch�T�½'�?���͖ǂ�k��F�˲B��ՠ�Ƀz8E �Ιlo��$ᏺ�t�6{�`����sˊe�e���3-� �3p�nW�!���}q�a�����A.�w%d(X8��m0;�H�\�أK"�g� �c����^�R��U]�y�����w،_�g~���D_J��r�?d,�C�"γ�d�+�X���vZ_�M��DG���~��3����3n��?�y�x����Ѱ����̶��,��H����vq�C�`W�.��#��$]�\w��nj��'�����(:�'w�$���BX��/&�2��9V��{cu(ݱ�a�Ē5���8��LV��F�Wm�u�/��Yٖ�@Ny2�~���l4�o���t�=(��t�d����0"�s�XS|�$
G�Ԧ�t�*��{R�z����2_�p�D�u��s6֤��?��ga��^@�<��`z%OA
��ע�
���O���v;Ac��O[�ݛR�C����#ǿD�����cE�jg�Fc�qg�0��Bɞ�@-�#@CK�V[�x��GEo��T�R�}XcG����c,�؇eٽ�epG2��=t�aȖ�nÙ�u
���b9mHQ�q~��Lʥ
���K2٥4ъ��5t�(:�[�=���@	�
�ҍ9���_^�p��z6}b2�)�Q�ΊVu�RdY���BfR'E�ޝ���N"+E�����E�G����z��3@N���n����NI�,��)[�{ģ�,��f�l1�I!�%�l_���Ae{wb�H	3k�bx�?�$��f����Y�M�w�-T*�`W� tY~/�dH�(�Ga�,ΛV]��٘�r�p�Ua�*>�>�&�����w�I�C��9=_�b�)����p8�1ɽ)���*X�#���c$o&_Ke-B�^ʄ�qP�v¦�|�|��Z+�|{cGq��cΤF��)���r@h!T�]�Z��D�)g��x2_о[_�vI}]x���7���k�f�({�=�rW���������6��V.��?�E�@
�4_��tlV	�as�mß
v��utQ�EO��5���j���g.��"Q�H��c��`�JҦ,�B����H�Yˡ�6a��e�X�@����b%y�#1���Z��Ц��-��Mwl�9�[P*�GǄ�_�z�"T���=�?�3�k:6O�	�t/I>���c�Z�<�}G���%p����ĠB.��8�|�z���g���+Q��7;������-TA[�%7��>�4��_���,����=�t6��zM�ޓ��͢Gf�\�\(���DM<S�"~*�E�-f���"����SU�E�����B�^�>��*�n���=�-�K�c���a�TF+	����T���'�e�Xl��R �aoZ�i� AƦ;�<��!��I(�L	�	����吕y���òӃ��v���f<����ez@���xO2�
����jk՞���l�G
s�VE]Ǡ,�%��!b��U�L�0��1& ��#&�n|��M�r^`��F�gnD����I����E4~�W
Wa*4�W��$>#������]k�9q��i�]���必*ٷ��s��+��J�2Ћ�}��van�[I�V/";j��A�S���1�H�xu�b�4��z�|0|߮X�?��k��t�7	�nQs���s:����%�IŮL�ܡjl�oA����6�h��*��<�� �}�e��6�S}��vot�ja�k*���gX.�q���%�j
Z���+j�wwу@�]��6tm����ȰPUM�~2>��s��:��c8��OV�����(G���O��|N;�(�k�������U"ef"2@{n
 �+�e%�g-����7�ЗH�@�x�N7�D�-��*}Ni}��1���]N�SN�Ս�d������(�C�c�[�b�O��R��n}�n�¸p���rYm�-�%�=@>���Fs�9�S���ǖ���v*`�==�E��<}<�����6�ʧ��&
9V�h��g�;~��� P7���L��)Ҟ]�u�6�r�����M��݁�R��e|�)5���w,	ֱ-ҁ���]��r�;��z��O��V�C�
�*�^	[//^鵤�5V5��2�i��Kt��	���O��׾��v�\˺�� E�x���U�?
��VPL�?��o�
*d1����q���O��m�`��@m�I�ÓX��ݩ�|sӒf�p�u����~x�h�+���M��cW�c�i{yF%�k��@���c�<��,��sr���v[?����´�����VS��S�/��oyW(���*E|��ĆhIT�,^w_GK�w��<�~���@�+���y~���,;n?u�@�0�lC�N��vQNj-l���n���\(i���$�0z�r���}�K)l�� 3J!�0��I[ 1��ޚv}%剜����7�c�tf�T#~vS��y_�Q <\��t9.�:�$SD9��P�R:�]�z�TKm�y ���}愯r��;�ġ�Ds>?��s���5性�Ț?k��PO�}���O_M��k)R��s�ߴ2DX
�M7"��u>AoH��l�29�:�#?,cu<X ���B5��8�c��q�=�d�>¾�{R$-�i:��-�#>d%��9ӳ_?n ��<�VV�ԫFG\��>_λ �kVϭ]�g�X��T����4�5�X�V|�@ᐫ��Z�z�g��;^��E>֪�tV߷�x([�����C�u�u�����'ǭOo�Ř(�6��*v���ſ�����ǅ����ߛY型��+,�[����XX����$�+��S���Vg�7$E�>U�>��
���Ŧ� �x�*-��Iw�2m�9��h�P�s�$��U��V"�9��X"���B��R�&�p�{���ߋ9�\�g[��/W^53�Q��x�Ā��05���&�/Ac2'�ʟa��p�n!]f9��$^�֍e�,�`�t�� ��k��PT��0�]��x�wL^�¢�Y�;�8�l���^�Q�f��Z+�ڝ��S#�Yl��qYh�a�0Y�4%���_�c$a��{��X-��m�e�P:�qy���svy��}S�R�����1j���.�� ��.:����?�ٯM�/����V�12_�k�=]��@�����_�[��;�e�^mc��y1D,^��4��=5�1p�P�q�`LIrVL��ٝ*�	Q��]����Ñjq�q
��˾�@+�po�����I�?$җ�A��0�8v�֘�m\���]�0L�w/�Un�AE�c��ڝ�%p*�w��:A�]�����֦�H��-�f�`L���߼O�Q���[̌�̅,vss��G9�;x{�hH�7]��n�$ɠd��t�8�/�&���	�pu�g�W�h#sm�fш�Å�L^�ɑ�:�1<B�h����6U�� c��4�O��"�rh��|���F3�W�.�;�I^�4O>M�H(�L�L1��*�Jn�O�{�8�!�)~��A�pX���4NA(kVjO��`�%���sf���P,*�H�ˀ-�u�gT���6���52i��V���ܵ쌜�[ie��2��HT3�O��D[�k��HhR���!�����"�P�Dw'�q"ɉ+�$�'R�L��=䎂J���Ó&v�"&�Ƴ��r�~�Tq���������8R�����<@�~��XE����D`6�r����ݣUEn�*9�Hű i�۔�5�'�v��s���� j�����KW)��xMQ�	HT]k�'�W��|퐿���g������)��� ���Dߝ�w������|O�8s�j�����f��(�<t���Y�MK��x~[*m�h���� �I���=�Z}�q��l�I��J��oB�CG�z^���MfYs��,��;s�]�^4��Y��q}�1�i0�a%]u2�l��G�q$�.�	���A��x�7��x������k�s�[�$�@��|�|�~{D��}&��J�}|�+���	�{/8��wsո����[�JEvD��m�6��h(jq�� ��De/+�u0>�f������]����� ƥG��Wp�7s�g�ډ��ް7W�m���T�8-A��L0��\E���Z��D*_�����B���J���Qp����޶6[MtlTr�^����C���}�	��*�8ع��*!��n���-�bCxg6f)ƯgB�-�:y�ͻ����|�bs��4^��00c�0�<el%�&�ft2��٥���9�D��}{��x��]LG �N��ҥ���!(��Nµp���iJ�>K�@��6�&F-6���7����.�1�ુ������~���*u^�<��G/�����lA|Pq���0{[����t�ק4�ji'8�5�h���ă���	��FO����:	L�Ր�~�ԧ!sथ,�-#��R����e\�]V������P�M��K`���/�������ö�'�^M y��h��'��~8 �4�Mm_��S��d�k!j{լ��� ��!l���c���b��BՙD�f
��aZ��޼;��K@�}�'*�r5
���� �֙���qܦl�Ҁ((�x���W��h���'���L4D�W�ʋ�v~"�
�����'�<�k+��9ƾW���G��t��K��ߋ#ǹw-�5c��R�����LF�Q���養���#TE�!Ƀ���gս?��&3�>'o:'�T�O*[o
�gJ�˘����42��s�N�'̽��XH 3R>��0g�Y�0-�P~L��k��j�7�7�`�GUW����6�Ϻ�,�O���fG�C��1���s�����6sqٰ�o����|1������f�����I��beS�'4�YS>�$?* ��ŃdP��R�T���XʛR\�M��O���0�"�����V�"�WȆr䞷AaRl�ڊf@�Q+�1UÖҷ}�*FsUM�§��LW���(ꢿ��"| >��:hL����;(YhU��W�-=��hW�`E�3�d"��B�e�p,��U�0P��&%��aA\0��i��Tۙ��&7������:%{G��A!܁����̣�쪥C�+�p�ӾD�&tSG+��d���N��i�yj4�?ە[�W�o�E����/�Zo}y��8��{Go�/&��pr�@���w��E1�<�Eb46�o<��FEY&��56�~@��>���4L��9y�G�{���,:5��݀$/������8�Ņ�Xkz��.�|�ƍ>���<SD��cn$� +0���=f���EEn�x�ȂT�Ӝׁ�) ���9�k�ip��n*��5L��s7B)�<��R�1b�tC�hY��f�!l��]�m_����B������?�I:&w�Sjs���!��&$kq�I:H��!#|3���e���?E��Fq5�2z�Gk��j��"��,�����QBS-c�r�Td�=$�o��nĻ-.�H`x8 ��M�ȇ����֩:+��/i��3�<���Sr���=��f7�8�涵c�B��})��UJ�C�X/�'1��D%���(�~�.�\�x��4n�7-5���pc��ǵų��J�:�y��M��e���N�y�&�-]܈��@s����s�Ć��\���������l�@�\�W7�7|�!��;��B*��DI��qn"�5��+�O�M�9k���7�p=�p��Ҧ�ɿ�A�X�(ʓ�Q3(���\��Tk���9�8v���%�&�+�SQj.�b>��.VM���x�����8�7�<���&����h����,�����+�-����Č%��ıi�N�� ff�= �WƉ}���v�:!.-i)�\�Kܿ��D<���y9��Y�C�^��5�pU;h���_�sj�0��GN�38���Z�"�P!�_pQ�]�},�թ՟k:��^tB�$������3�k�)s�.@M��hg�zճ hD�A�~7�qH$1s�J�x�"OHvlv�� )F�3�Y(���TJ_�Ty^��`p�S��{ʌ�m�s��pg��IT�O�M��J��Za���4�{ů�شs�pj��;���E$� q8��"�7�C$�׃�lN���{$�l\�6�����yÈ^�|�L��y��}�y�jl��y�
l�lh�d��u�{\��!9�0{s�nۻ�HG
�rd�]+�k�t��?!ww��8�� �x�~�qǐ���'�{��0�UE�#���s����"���`4@��$t'p/����K_�f�{��'���cI=�(y'����J������𿤼e�e��*���l���߹0D�7+�¹�i9E o���Zؼ�C~�ru�Uõ��u���j���l96:%.wgE��w&MV��?�x�bAx�z�Y����)��@�=�榏������έ���DO�<�D����b�㼾E�OKu�-V�Rb�}D�@eH�;K�4��&-c�������n&��@w���[�7R߲ ��ʼX�fUA|PM=��W�Ŷ
��O�G�K�j���G@��X'�.'�XN�r��6ҙ+<��%&eA�4�W�v�3 J�ǣ��Iso�:�C��{�Bo*{��C폐��O>���)�W,�?S<�<!t$�?�����)�͟􂏂������R8p���1����E�ZbXR�t��;�x���4`I/�UޫJ�k7����n�|��/������M�|��_�Mi�'rł�y	tv�>yS�}����c�l��z�#����G������G���t,��~��*����s�l�'<���?�r= V\�\	��|��j�$�	�ҙ��p�:�#5��Ꚃ9��՘�B��J�Gi�z�~,��n��Îrք� .��a�0'��8g)S\]�h��Y�wp}�4���W�T /�-z̗n�+�}o������_�/��J2��Ԏ^���9��mZ����]���,h��Z�!�`.�ՠ#d�	ӌ�����a�`�F��R�^g&�;����yejiB�1�F�G��� �0Yp��bV�(�(S��NR݋>]C�V�n����B���~;2����v��lz�����%���Q�Iz�l�}�`�ڑ���I�Odqǚ��K�W�N�X�*f}j��V�2'z7��w E��R� %�>�q����9���˷��;{��ߨ�B4J�-xu�J�
Bogޱl%����|
�^D�a#w	��hQV�@��"D�_6ܾ+S?j,JY#�-�����߇��fP��Ü|�`�'kw��.j��1�X�)-BX=�ɑ�0�3�b�
^��� ����pӂ�	���e[�3�`%��<s�:�2Y>�К+�B5�N�\�#	v]�EP��[Y�s�v��;·�����3��_؇'�t�aV �n���f�o�P��8�`�ץ��b�-�+8A�-#n g�1O�ax�է��**�8�ڕ�í5K��j�=�?�Dy��Ɩ�7@��J�X����<	�
���i�[S ��������xA��N�w��;@��������8����d\sQ��x�C��'��>� WF�
c6�Rኇ_h�ŸuD!&����� �x��N:(�3�۝�>�eU[LH�V:���~Y�&o�.��ܘ[W��^��__;W+#��-�Ce jc���Ow^�!>�c�ά���Ʒq�LCL���8��ow.m�0��
�F�*@�ӧ�9�����!*V�xe0&��&\REV�1v�3O�	ri\s��=X��e<��Ԓ�M4B���(\n{ޖ��3aoG]qȎ�d�fP������j	���y���C���do��:�3���b
�w6�ܮW4S�=�Ӑ�fyG�ƪT~$~�Y�k�����Dy#�ˠ�ջ��*9��.�/W���*b�#�5(SM�-Ֆ\%�3�?f����d��xgc��v�{z(��$�n�t�Cbv���VXe�ҍ�d�)�$`3�s�k�����(��j$�g:U���VN
Z��[<�jg @)��jh��SqW� ��z�����B.(E)r�x��1�ʛ�)�9���8�(�1��7a�!5la�Y[ωB(@�{�w����/�*�SD�8��fy�!��$����ṬT�k���zX܄��n�5;p(�������>�r��n�0�H(u�H��$er$(Αy��.U)L��u4Q<��O|
��=Z��C�^<i��c�Ky�m]lm��D���v�@�=¶�r��,-�Roݛ�(L�>4�G�p�-����-:�/�Cw��f=�s�����{�T]�z~�@�{�t�h>9yI����
��T-g�3��>u�+;^aY��"�?N'��0��lūo����n��ף�ū�Kqyl}�N���������B��R�/�"�B�?��2<�˂��U#m\�J�����;��tX��_�T�v=(�����I���D�C�46��Qr�4l��y{��}� ��s�����B >�~��U�a��kS��)��b-22#ތ�y��o���L�Dz����ۛE`��]�u�8~��{��X��|0�y�1��┙D
c���©�~��� �b�3y�I=3�a��(��k��E]6r�cѨ|�aN�Jn��3N���m`�A�ƥ�=� ,l�ŹZ*��Q��%y[[V����,�T��"���?����J��:M�������ȝ�؈���x�F/�m��. ��5�?����r��J'K�uRiB�e#Z�����W����do3(��nm�4��J%���V�&,EJd|���I�4�{�d��&ޮ=��*�uI��UR���8)��q�?�uԫ���h&X���Kq������B9��M��!���rR˒Ӳ:�|�%���_�D��uX�_�ir`����ZHF���J��ln��7��f�@���~p�c�5�y�v��̈e�Vq�J�3��Y�:Yap�&e��-P�^��jD�ؚ��M#B�����|`oFz�]+��	��Ȼ�� k��K+�m n,ϏX��b�8o����ZBʫ�D�eB������FL'Ǌ�V�ͩ�|��b�h��^���%$W����lWld>m���; ��U_�+
 rn���A����F�iJTl��1��"E�o�n4Y �F�/L��g���2$��@FΉ�m�MPg����X�M�P(��+��j�U>��^�n
K61� 3Jo�Z��I}�h�J`S���d ��M�6�6��ҒA]���e�wsrXn�}A#t��R���3\D�����&�wS�ͩ����r��zR�����PSv~d����ݢ�K�s0V����[9^T'Y�-�\�g���e����M_���?����6�h�t=�-����b3�|L(�9Ɖާl�vB��y� �]"�=��ϣ�����
sY�A��!��*Y7�GX�b���x�W]�&�+=M>�@P$~Y��Am9�@b��`�ˍI�h�Vou��@�Ư�*ݲ
���<DB7�}�V�a�\�..G����fU}���~�ִ��$c$O�������0=�op��o��>U� c����HU���k��="�AF*?��qt ������
( 7�[[F�$���x��N��
� g0��K�[�_�Ŧ��SG �n/�:B�W����P7���*�4!���c�F ]�v�����-�Ba�� ቾ���|)�����9>V0���	��k�Q�dy:gU�n�\��[E���=H��'�#�@�i>� �`=�_��%�M�	)�*����Sc9�5�|e2��cY�[�e�*�X� ԡ���P��� ��������Y
���h?Iu1��d�$��V<�t����#h���dPb��Jn�p�ƉB�aw)�h���� B��o��#��"0��T���.^_��tЍ)�*��^f[9ż���V����/X����*���LX�`zJ2��y����c�Du���6#r�t֗������G�p��+��V�Kȡ{�/�GP����4����j$���V 
9��,�B��������������%
g~� Mnq����#��{׉&i:�ѩ#��Z�βS�؀UO#����ʑD֛/���Ϋ�I�.q��� Wbe�+\������L��,�ۗZ�Mv�(b���	��5�p�{�}H���Ze��q7�o$��H�5K�w�X�9?���;qI�4�w��y��<D0DRaߨlnc'�������U�&��2�~��^�����j�������)JH��P����-���w��K�|,���A�"�g(�_�l���ߍt$qU���^�}��QH]�bS��l���-n�Aw�A�<�}�%>˽�8|A���#��Ke�Ц���3�6"	Z���qP�"Ο���a��ŧ��o�	�>��A24�ٙ�U��«�_s�L�aK0;˕�h�,j3{�Ƶr��:pց"�d��Fǁ+Y�st�.���Q Yʡ���r[��w�x%:��66���� �i�F{��Q�ڋZ��!'�+��d(�.���2x�����N4�ϥ�D;�A�X;�$ .J�]��#L�|���X�_;����t,}u��j�S���1o�'�(��]ʌ�Eߤض=���PK"��$D�y��=��~��D0+��qV6�"�,�z�aq���5Q>�2��t��B�O?_{=�梹�H�Ъ�Hg�BXG�/-�H�mmæ�W��n7��+����d��}�v*,��'@UB��E��?0M^r���%�?x�J9!'��w*�ě� �!��M������:
x!��,Z���a�22�q57HE·�[WQ򆿂��|�rX<t��D�;��	N�#�Q��ݪ���薄�6tAA�J\V��<{抨���(��\��0|dե$6'J<P&,�\5`cqǯ���<;ڱ4��/.��A�ږ���61��J�q��;1U�o��HF�&���SRW��G�:k��j���M��e��N���L�lh0����wP7��КL|G%�J���#`h�+��� �� Z#s��_htB0�oߍ�U�$��|���N]����3�\e��d�C��e�l��% Ro��l��7]-N�:9w�1��e.���,;i�9�Ef<�Y�s�`�}��D;���A�:ؕd i�x����b����������Ḣ?+�iU�8I��X�t�O�Ah�1�52\�3���]��3y�ncmk�����o4_� b�\���k0�}��&z#�K��]n;�2�?$;X�,�P:=��9�P9�4���㻋��W]�8��0�u�w��~5g�՝���:V]E���|�Vd�*�F�ѧ	�~|�	঎'1������!��2�����J�	:L��i�`$s(�CvR���4<�ַ����  �w���=$�d��T
�UL�P��9*~?��Kv­�\B�[��\��8�|�)��%*@ ��>����㩎�3V	�#��3�d=�|=E��k;�������'B� �?ɛe�֙Z��ֱ�����\i��wֽ�>�V4�/���H�W #��ttk��J�^��))"�W��?�.����]��3f�9:�Cdy6���̯��g�]u��@�+Ux�7�����m�ʸ�_f�{	�0��'��"��)�F�ةI������b��_'n�by�x���e}�=�t��*c�{��0�R�i����czԍ��g�փzp��77(,�@��Li��M��/��J��P|�.�|H������Z-{��۵!*�F���林�/�&�pu�4��p�W���^�����?yQ12�Ν�oz�J�+�!��f�6?�nP~��+���g��&m+��I���{g�@i)�)��A��|X��t�p�т���i_y`!����K����ӫYe<�?g��cȕ��ȇN�m��ՓX*r�G�+��K-�ݪ��^�w@P�m{ r5L�֝�zjo��O؋m��U�>P����v���j���:,]��ց�z��<+6�wz�����tܟs�'Όlv{�J�8�D�+�I�4n�����[�f���>��6|��̴Ү5���%��}�V9�g�}���<�3���Y�0+kV�� �*�P�������z��$���*����������rL���3����܅���i��7�bS��������Z���e�8�����D�g�+�L��F.�N{H�S[�<��RB7�OIC��A�>�m�%ߋrrq��	�[nO���W��⃢����x��)A7�}p��>@\
���JsD n�Y�kN�~�]�h����-��ŭ����թ��!(MV^33�#֨����g�ِ9(ֽ���2�w^J�r��2�Ru5�c�w��؇�%1�z�i*�@ݻ:WF�ڿ���M��I=)q�T-�������������*�(<��x/��J)���Hz)GUJ�.�Kj[	��Y�;�3[Gk���}]4�$�+�h�]p���}e.��A�� U�5r,�N�C��HҹWC��!�qyWu��C���e���Ձ�����'h�<��~�e�{*���cvR��y0N�Mf��֑�g`u��$~"f#~�y$��)8�ɀ.�&^|���ٿ-( ����8�p�����h���lɋX���!���pM쭘]>�� ��h�
�da(&C�ר�e��q1�����zf��y/���f2�#�.Bi�Y=DY�`L?\�<��+��W�$��)�&���-}�Ө��(�[��� �-G�F{��H��߂�����9�$��ӯ��q�`v��'���4�,������{���'�`�l
-z��U��(��Ҝ��2�`M\����@%n�޲�)9�#���I����B�z<J�j'�F��)82G��� M�t���?�o|�Ju4��L2B>G>�䳪��ϒ�G]ȾΗ?�!�9�ٝ�k�e��b��%6�#.��U�kB3Q"�X�װ�~�^¾�zuk����4���FͰ`��Y��4�|��ʝ/0�d���o��}�aNkr�&cN8��'��ڧ[ۜ �s�wIu=�W�z����016�I�n��xUAoCT�е�f�X[�+�%������蠖�t����k��n[w�)%��ΰ���?RDxW�ʆib$�p���g�S�3�oE�pK��<�� ��'���B�� '���8�;��7%�㹆�k�L��	�e�=8E��B�����@�%�΃j��̣ow�M[Y��I|�Nr��o�N��o��@��T�p&br��{�F�p9DꖲO<;̹�߇�/t�B��p>V��&�)�L���oIm!��B��ˌ�fA:_�[��)p��+^V ~Ur��Bz���F�\�S��%�@�T�#B��r�.�@������@<c���WD�4"�ܲE�t� k_�% ���x0x��I���ׅ�1��!O���y��&���J���)4w%G���V�"�*�\�Y+�iOź�n���}D�h<��n��9���6G  'ͼ:�BٲЊ>hq����!z�Bo����B�α�wZ��������ͬM7,�W�L)�1���B[s��I����b�9��i�w���p����	�}����-�Ku�'Nhx�=�0��������4�
~^�$�hg��N���^���{�B��N�5�q��J�Ifo��W�g ��܆/��`j���/qH���e6��Q�����a�OS�ΡϹr;!(n��$M�H	�Bַ��쪂��?~7*'0�J@j"/�W���4��L'q�7{�^�L�!L��pz����
D�Q_7����d�K�{�4YZ��;�7{g�#܆�3qxs/��*p�-r��b.B _a�5��aP���b5bpZTT2 M�|qڱ�oa^�����Y?/�'pd�d�b�r����/Ӵ�6!m!��/�)�d^[ �+jq�~�C��k5� tm�MTVGf	: �ؑR�}�a��3@RFԺl(��DY,&r��	w�>Ld@�2*p�os���ǰ�{�ϝ���Y����.�����������b���(W|��$�Tx!W} Q��H?ғ�|�M�2.��h�=T֐K%okM}rYf�$���L"��wj�a�-�Ɓ�y��u@�����fI�¤�PVo��}�^��F憐W�hj=#�mB)����v���c�A���V���U
���A��K�k]h-Aդ���	#Z�~�h�R)T���H��H�걩�)��C��o�4��[��B���Z�� !$�2yQ~>�"Π�笗�a����o���ڭXQ`�B�-�����S��*g�o*��n�����Ŏ����S -Ww~��L��s+~��+^Ml���gN6�eAC���On�h��}�ng�!r9�IU.���y1s����p�9g�lK^1{�C4���Q��2�I�&Uj%!��V+%�Nli# P��|uj����+��p���Vc.?�֠V7�'.���^˹t��:�`��Ee���[��<.d��Vޞ����{��i�������īq9�_�5)��8��� �ay�3��b�8�}�:����*�t/n����㍗�f�7��^�z�q�
��v��E���g&��x��_�:Be�eFG<��]��P˸��:�o޵CS����f��c�Y�+��۳�̊�Oc�P����:��K��-�[�g��+�s�T����	˔����\�B��	��W�(k�'%���'����9?u���0�3���	&��ͪ3c�`��ǎO�u{�Ki�肳&��q�[(�Zck[1��j�3%�čf-��~��\q��S�rʸ���'����B@|X! ���^AA�;L��ln��4����>�W�� AJ�f��I�=�G5�p]��:�0/*j\@��m�&\�tm+�q}T9��kh�1��]�B�u��Wzĭ+$�\H8��Fi4�C'��	`g�0|'��ngk�$���ا�4p�,�CI���@��+�_��>���Q�;�<�cß�W�R�i_� ��:����XCHF���en��tF�uV�~xs��x��H �G"���W"h2WB���AxK!{��a{k~��5�k��G	��i���q�Y|a��9@:7-L�74�o���^�1�Y�B��<Y -�+6������B�'A�ֆ�+{��m"d<��=�Z��YO���f�Lr3ؤ�*ǐ?t5�m^M���{z�:o �*�]U�q��pM��v}�BA��#���sＢX��=u�S��R�a|�ϴ��*�v�M���.#m�n>�ʺ<%�C/YJ���3g�R{<�������.hjk,7B�*��=8��&�L����O7���`2ה�������\>�|��sF_R��aH��	dKj,ɴQn��H[q���j�_��Y6���9�;]���Zv|wA�5��WX�f��*?����H-�}��b2�6_by/dJN�������"ߟ2�u��TX���_9�����Ͳ^�(�a
'��)�z,������S\kF$�� ��W�>����j@J�)x��rR�ǛPS�^�ɉٝH���-H�����&��zu	%����#�nF^9ܹo	Ɏ"�%��}�N:�o�3Zv�=[��*>n�!�~��r_[[�8�O��q#0(����e'v��U-9a=_a���c|��$ƢPK����T��_�t�P$59��w{����N��%�mP�T�k�2�K�k�M��E�$��_��]K��[i$vV.��_������C���F��3����}h�O-����UQ���R�d��%�`ю|{`
m���$f�f���j=T���@�q���a� �p-��JCB$�~0t�Z�<�&���dV�q��}������\�9`HP��h�3���_)b%I�p��?� ��p%���ݤ�$���{s"ԟ�s.5���eH�oR��v��F�(��|���ۘv�P�3	ߓ4�{�:�����=��vI��r�^������i�	�kg?19ۘ7EQ����o<�D���编�
�<�r�",�tլ12��=�����7�]�����9$Ԅ�2lrOVMc	H?S�Jh$^!���@,s��;w�����/���P��Z��7NlU��A�m���Ƶ�9�Hy���0 ��%��X�^	���K�h�u)���jT���8O��9L�W�\����Zp~��O+�����&��4�>��"�F�U����6�k����`�����K���<O`ː�\�kg���tg�����X�1�o��q��x4T�	y-j��
w�4ͩ�K��o"�q)sҟ��������F-p�V�6�IG҈�iWd��1y[]�E,�7n�����}��D��}��a���T܃w�~=�'O�n�>��U_�Q�6/72w�v�<��̅�6�4��W�n��^0���f����O!�_�=�gk����8sqs�aU�ܾ�ףa��TM�	&�
@��=d (�,�m�
�
 ���ru�����H<�j��כE8Յ����J��(�s��[��>CavB����p�=�I9�(^g��L�Q��8RO�ܤX聋��d\o9%!���� ������M�
T|3��DiqUKt�q�i�Z1�%���p��13n��>��)�=eA����.�&���	-�P5D�;w�ɟCJ� 4�*��tq�)�����P���>e���V:
u��r���<`���NF�!�R�%��d5���F�����?M�Y�Ūj��~���] �/ZJ.���o4�{sיɪf�r�폭p�.�n��W�k��HnX�D~-�q����"7�D��V�P�y|6��8���.-;��A�`X6w�EVL��R~@숓v���%���q0�nb�Yܭ�J�OU��"4l�ɱsN
�"�^�x0��1?��Q���FW"���C�ª��!�T2>�_ߐ��C/?ÕU�T"9:Nn�7�`�Ou��gwIƊ�1�1��S�DD\8��Qou�HX9.��ab�ot�yK�� ,��C��cc�(����J��C��;��?���i�.��W�E���|����~��#�	�]����A�ZP�b(�F ���/aq�Z*�8R7��^'�-���z�=�\�%��T/�0��Z7j䄆밟z��I�1�1Z�/��x�zw��Vy�ƢS;u�����������/�����>�:o^n��;С��?9l{}ş��&��Z�Ϭ1�I:�Z�R���B�BS}p��\Y�V����i����,PIMz�L��q��"�a;�\^r  �����e��V�&�%|V]�K1/��ͻ�ʨG��H���H�T��:��\Rb�˔�����C�T�}s`{�$\l�6��X
���Wˋ�ո>�·������E����5e�j�g.���m����*�lm���V����J`��G,���7d�f�O82Q}bJs.��y�+�u�<��5�w�f|�>	\��Le�`� ���ۈ��LN�C��s�# ��9?v�H�э�>�?֒�N�;��%��idL�)��z?��
�!C����������2x��(3[�E���j���]r< U�l�ؕG�{�/�n�n��F�oU��G������e���dF�_��n�Ee�r���Z(����s��~#k	�8,|��W_ܢP|?��j��LX����s�����%�_aR�rbX���|/���r�k�"ز�l+p�x��t��/�~ao������W{*���jVJ����HoL���&�	����lq\8;��-��vwzBWiKu�������H�R9i���Oÿ=�\�И�~��q����X�z�ᳮ�ti9sY	J�W���9�O�Ici���-�d������ݩs�S���[l�>�i�ը}+hL��>�G Alg�ޚ�5nKg���tP��,�py�8R�]�������Z���jׂV�h�_��������=�Au4�_8��бײ��۵�K���g@5��N�@if�T����A���D�z��FeeI��@�pF�WF�W��Ʃ���֬������P ��_/VO a�h�<N=�f)��Qlk*�[�����sG�b�>(�r�<%O3'����������hz�
-�i�"z�pl4>��_elL}@������Դ���ů[�dɳW��?�#)�6�"&i7�/�TfOe�D)��f�|[�S�U�;4qGL}��fǹQ��9�渠�'Wp��S5�������.:_k9�����-
0y�ъ1�4ʾ�}�����w��]���C%vh?�����|҆�E�q�3�_�0|�rr�
��H���W6s��4r����дH«R� wWf���0�;Oѵ���5�ɨ�֖��m�7�9�{&��Rs���$E�����uc��/��^�eNg�=�qр�	�r���7�Ҝ�Z�C�oS����(�	$6W���}Ğ=�*��8�%k>.~�{���h ����V5���4W�� ��4���?F�NJ]?��4Yk��� a�E.Ol�d�x���qP髐U�Y�>	գ��J�+��(��)���Lo9��� 	��;GOexٸ�cV������w��G�O3�b(7�
ɒ���B~`�M����sI�!L�NB0>��f��|��`	��4󤰦i�,Z<s�ti5n�Bl�ՙz$�`="�7�7WO0-sU}=����h���I{��9�l����O��#\�J��MI�&�^�~ҦU��_V�ux��Ŵ��޵taaU�SN��RcQ}ϡ�l�J�6qJ��-�R5��>�ك6�e�7����PB$~��L�I�Sk�Y��B�Rd�$P�)�ԝ�7�[����&R�pc�3��qZ�0!�r�O�l���%|�+NM�pLi�j��0&�G�+[�4QO�>��J�,C�h/��m�#�f�FZ��vk<ѿB?��Y�H��^k����P�I}t�Z����Pɮ@���-W�Ô�J�8�����FK�z�w�O
��'"H��ܞ�ơ$�a��J:�`C�;^�8k6�x���G7��KI�-����B�N}�@O�-���[+��!n:����.Q/t:R�ko>v
�:y��;~�q�,FS!$��>G�
�G���w��ƫ��>@�(cVZ�y��⚸���8{�G�����7����L�`E����d�	'D�0�_qj�K�H�R=�Х�ȥ�ϭ�^_����NM�1��OR٤9�U.$�V?RQMu���������e���x�V�(���׭�E�@q)��R>_\�)9f�q��5�I������	gE�B����[�r]�*�R�a�^��=@۹��*�\�w2\D��e���x�#zK�/oHY��-�x��������B��c��q6ñ��TJNN�S��%q�;��I��П��l�A^�s�u9��g����4����8 �����1��ĚVB�]h>)�����	�EH\���(���J���B�Uc�ZM˿S�#��8ǉ�������S�����A�m8w�K�'��;�sb3W�?��~� �Z{�n5�UA!����},������O�=��R�?3���w�U�H������r����)'.�#2/T�pj7�4Ljc&��2��}�R�8>%�;��Y�_�����?u�_�B�A"��=`���3]�L8��N�OWUV`�IcT;L�|�:2�@R�e�wi6�>oRH�F6�����U�N�����~����ԧ��"HA,K+ѻ�mk?	x��g����C���TK�7�0��?�sdׯ+��ˏ2��=����h�pf%�W<�L�ob �h�k�'W�<��=po0-P3��x���c�2��>���p�Q�T���r��baG^?U�<��t��p%� 4Q����~�O0c��мNy�����c�e��.�yS�Vd�,�MpDn�NU�l�,D�_�rw��}�z�����i̫�ţ]PF%u��}����6|m,�?],*�����֎�V�k
Q��"��і�}_�f�c�x<�<��I�!���<T��[�XX�5d�ڂ�i�8(�S69���+���];��C��F_��Î���Uk&�8��|Į��c�-a:��S+�]?�)��sO��2=�;&r(Z�U���F�_�B5���=gtQ�B����=-�k4GcJQ�g��JM)1,���t@�� �aX�t��j��}�X�X����3��*!�5��C�mI�i�4�����0w*���A���i`W,�V�qL?�Z����ת^�Ly� h("��X���!�q���v_o�h=�8\�������B4r*�5����o~�=�B�Z����{Kr��s�p�e��h�L�7��~tx�{�W=cE�*\��<�苛�kuy>�Ԍ�_0��1)��d~�c��^�Ip+B�si�~o%���4a�)m��� m�"�����B���S:Ƃ'�!ٖ̙����:���������v#���z�.��V��G�����q�Ȟ�����$����{8���2���Yl��eȻ�V�+��Z�x*ŀZ5�����:�=5�,l1}.�>,t0��r�E�\��4�i�]�#8D����v�%� &6�i����wtW=5��U^Z���X�R�5P�A��&3��e����ppr8N��i!z�5�(ބ����P��U!�~�����ޥ�^�Ƅ��d	g�\]�U�+^V\6�J�b��jZ�R5W�����
�f����c�C�B����b�9X�Tqk�rA� w8�/�����m�{�����©=���ɯ���K���&�a!��5㺽~�I�m�e�(���i!��S���y#Q�u:�[堄>��4qq�ufc�fpتW���b���3�MG���'j\�w��>��4?�2u�`��	�G^����K�$�ENYL�B���TCp�`�"ţ&xt���=$%�z��x�.PL����]��.0�~%*/��qK-}8�R����a˫��&l269 l�ʓW*Y�l�e ;~�K˚-'�R�x.��Zϧ��f@��&К/ʻA��=�^����Em*�4[���WE�"2�=��(��jX'A��q��0�۽���������xՙ�>��8�� �=K� E$�w�&��|f���0t��#��6�_�+��	[/�N=6���?�G�<���6�3o�J��h��U�r��w�����\)�U領�<
�>0��a�J�����J"�6�d�	�7�p����m��\><�L���]�6`_�M&,�;��^\�O��l���!�v�"�WI�(r'�%U?_j@V#���Ɏ�G��%�y$M~y��t�Hΐ�;�y��ZS�dZ��p��j%Rc��e��<�|B����p_l^{OH��
a�q�t���^����d'��w�=�Ԣ�~4�*�D}�@�s�[)Z��4�ԣ�6~����؀̈́�	l�5��f>�p-nX쑄J���޾�Qhۄ��_��"��KE�zD/z��C�����y�O< 
I��G�]p+Ol��?�x�<���Dg@|����,53#�#���7��3����!���#��!	���[�!B(X{]V>e�f%7Y���n��&�'�o��p�kJ�Tr=�X�T��/T$���n@w��9Nn=,�а�26��"�r�Ty�B+;�e\d=b�������e��ϴ�V@<��,:��4�{��6Rj"`Q$HJ�n(���\��^�����@>���%a����8�<��hS������1����^Qg�ἥ�`�(v�o� ���[�dB֑ȶ��I#�K�ߏ��qw�� �V���ŗ���L�&&�kY>H��N�G�ꎚ$c�F?��6��=�2���� 5�{���xi�K9��N�� �o�?yay��ɢR��1�mB���{v��X�WT�Y�3SK&(kO$�ܨ�o��z�e�{����3u�\D\H��ۙd���B"���U��e�����I��n%�Ͷ�s1����,.H���IDF���Z ƭp<�������,ԢS�sJ�I:�)�P�>]�@2�0#L7?@�J,J#]}���[�]�B֑��e���3�H�wqC-{��>�93�3��c�wWB�o&��} ���2����j�F3�HY01;��Ũ70����{I�PÆ�?0.�F��G�s�[�;�x���5�r��������eD���ՃٜR|qЕ)Qd4�e�� 8Ԣb��] �����E��%D��S1`�kP�%�������-�/�lv�<��D`i
���#��G/�9_ז:;�t;he
��m�h3�|��{���N���}�&/�0�q�.�Z�'���>��T�Z �������"e�|hdV��	GpѩM��ݼ��Cٙ�Ϲ=����Bv�%2]� ��<���5l/��µe��q�w�V��~���c���Z��'y:k�q'{��*�d[
�N�ծp#%n���D�0�0�	������i^�IVЗ[�H� e &��h	Z8��gi��W�lZ��f)�9#�V��Y��0kE[��B�z���|n��駹U(q�q�S��c�EH��:��ܟg��fy����0����(��[�X�]j��w0�|M�7��T �yƤ��J<5j��)y��E(Ć�:����~�l��A�=&2�ǬO%����~Ůꈹq[i�[�����T{�i���������z ����\�]�l۰Z�GW4��-����`{�$���QT����s�I3 �vU�$��Wδ	��s�@�ֺ�T�R��F�z� ��m6�m���p�=g����<���I�!.���Q�B���>�7 ��F�V L����^&���� ��ŬK�m�Ⳋ#)���I���w�Y+H��Umc����(�O�A�`�O�k�p-c)6P���­�o�����2���N�r!7�zv2�e�0��U�8b��|��%���B{˞R�ؒ'\�_��0�����p�:��FфS�b�.�uY=�����S�GqI��7\"` �fʻ�.
Ѧu�:~�xwc��E�z<}���kz�r�G��O$��R	�f�1�R�z����I�l�%MGZg�:9�{�a��G�Y�@���ǳ��*�*�]
�i�͜�s�	��S0���D�a��4{����5H�P�z{B`�.�_1��y�=^1	��V�- >��Kr?�W/h�l��J*Yѻ^��u�ɮ&YL�B��������f�1�v��8�����$(P�ո���ʦ+�o������L�NL�������%2��O��&��� ��tL�$�F@ͱ�
�����u��7&�&�t����ju]���U=��S���+s`�$>��7�h�
�V����j��+I��6�[j���$q�b~�3<3w�7�/��(�>��c�M�~ۢs�X}9��Q���(:�m�qY���t�'WS8�	K�:e�j��/�6A�auBq>Y76b�q`�L$�M����b2R1�6_�K�bf�A��v�������c[��Նt��9�뗛VL�����Nj��7��h��t�v�	0�]���(�S$��S��]��a����o,cS{�!Ӫi�đ0(����Ts���X�ҝ/��tH
�E|E��f,Pߤ Yl�·�����݉����d�
��W���!6#Ep8K=-�G���%���!μL���tK%��/�r���B�_֡����ޗ:F*�z6?�3�!!�S���pw����V*H�1�\=�W�n��]��D�y���bZ�I�MM ��C-����O-<���B�g��X$C#6U��+����X���·m!}�+[�zӝqX�i���~��X�������=`T��?r���t>��R�
�50�v��
u�9��СA��۶^���+zL�r6���꣚	Q"���4U۞�-�<�*�߰b_��%F���JU�DZ-��Szl�����&�┮�q�Kb5�!�����#�lUԁ��lqI�$&��&��,)(7���r^�NK[$h���/<�c����b��Vl�YY(@5Lf��;�b��/�M-�y6[B޼��
���[Oh��ǳ�������w����ymA����B��i:Z��k�o�q%�l��.�d�܎�U��<�|�xt�t;�ZC$�1��Veg�Y�8�[��޲��];k�h���"�i ,:H31(��Jo+�1��P��E����de�/����W�0@mͰtd�87:~�I�;k7��ʺF��u"18y�!O�aV��q�[�=Z����|���� ���܍�񘹑������<�;�w{��ْ�g���]�l�p�5&�MBvĖ���n>��'��rմ�8�Ҟ#�##��S��R��ID?��+j��r�D��@��+X==�	�"O_�}�b����G$��G���-�� �?͓x��2.5Ki�V`=�v]���jwY�%� ����_�;c�r���A��TGo���`�S"S���t_�ˏ)A��ʀ�.�8	C�K`D�\��� �8M���#5޺�@�ԃ�,��)��жR�y�&\�{�8Z�=�_�CҗU���N-�	01i�c�Ή����y<D��,��K����>��Sv�=JAޥ=U����Cg��������W�ӳ���^*4��&a��Ŀ3Wf:��
�v)��)�
*�8��/�O����j���8�On<�[Bc�:��D^;A{Yo.$;����6�btO�\F���j�|hg���#"6�.���z�J9k�w�@w�:	�TŴ��~��� �"+��Hr	���z;��q����BWl�����7��[@n%A%���2M���`���O��l��A��:��^o�̥1��?Jx�f�j)E0�r��*���Y�d��K�.�8V�����9z�Qä��3��c��/X�6H�E�m�	E�p�߬��?҉�Aٸ!�u=�Z�4�����YGh7[t���q��tHƠy�c�O`C�A`����P��PԐ;	���Nٔ�Ju����mJ37�}��gi��!`�k(�-�ZD�r������-8�J[�?P��G�����(����`�"�H�=�妵i
�6�H��1�Y��˹m!�cc�1-��ވ1��=�v�v�[1t�m����E�"뗧?+V�����X�?�i��oҝI$|f��	�u�&�$W�����a��ۍ��\�&�N���F�gg�
l' Ɛz徫7�xr�m2kV�-1����;l&4EʅA4u�^ʃ'+$5&H5T�b�>ǹ5ag�x�s��Y�Y_�t��?N����̉X�3Ә�|#v�~G�o"T����Y���ʴK���ԣh�1}��n>6b�2h|�0R����$gV՘��Jޥ�|�]C `he�-���� �u�.e+�e
����UM�A}�k�ֹ���9&8`�&��`՟�"�����m��4z�2��A�N�K���G�Z��{�����Lš���k���@t�:��@k�񭵑��g�Wӛ�[|�>�Y��T�T\�OP�E��X��A����9Mb��BN� 6������ȅ�=su{.
ysx�|J�J�]S�Jw	1����D;���\q�\���(��T#, C52�igZؘIa�X:z�������$��q\��T�r!BuۣU���\�z����ie���l<���0���;F��'���3�W�	(;��l�re!�c6۞���?�f�<N�k���ћ�[
��XZ��W	�"WY��`2��x'�µ�����y_Җ_�x�5��Xs�|��v�_Sَ�KX�?�p��C��}�Y:bK�E������H,�2df�� ��)?�N�\��²/��R��!��$�(�;u�G�c5������_�����P��iUҿ#j��l��LX8�#�o����������aV�9��=�|�s�!�d��1�{����9�T��H����#6���{�*Z��M�S�ߠ��-#�p/ҁ%%Fit��92��`7��I��t�D��I���n$;�N�A�A�l�,�e��9.5{��|�5V��{R���`�]��=g��q��ΐ����V�aqV�;:p!N�|~xP���W#�,Јp&�*`c��T�*��@ٷA�9@��d2Ƒ�{�?�J�s �M�W#�R��Y���[K�p�u��7e��������c"��>'�S^�