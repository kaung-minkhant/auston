��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%��^6&���z��R�f���5*�< �1[J9���!1����!F��x�*���x�����l��}�:���<�<�k�)���n(�7��*H�v�Ug�+g}��D���(�<�Z�1*=�}��)�ߕ2�<��О����۝�f_�s�qВ�pD�:U���Z�.��)�x,�tՠ���Ʉ�*뻞VG(���Ļ���iH���W"�}�1'�^����͟�襐���9�1�'k�V��n����}_�Gե8	}P
��7&��Uk�LL��{�y-��TC�lE)�t���O:|7�m
 q6k*�ul
N&ρ�r��T�j_t�6�a/z�vO>k.��A��cMGaY\��6Pǚ�0fT"��$9kR����`P�M!E�S)v�x6縳��7��T�[3s�=��}m��Χ_��-���=���b���2�ٞ;�!��&l���A��ݞ��yO�yB�2{i�h%���]��s.��2
�*��e��y�?U��S�w��>������)�K�p1L���[Ŀ^7r${*�~t�f5c�&�7	Yy�*ˋh$���'�J�ET�1���4v?s�<}���l�lº����yY��~\X��D˧���T�T���Ґ������\5��S���g9��5/$@h�9��o/��4�.�3O�^$(j}ѣ	d�ž�㊤��j�io�������Dɓ�m�Khy��F�C�΋�%��s����vCC[���H&��Æ��hg����^�[�v��T���6�p2��(������(���=�}�җ�Mk=�+㭩hX(7��C����[do.6͖��$c5�2ƅ�A,]����*g�.v��Y�?���4��HXNjZ�a���N�>����7gF�G6�!��
��%Y l�׾�NX�0A�J5�02ye3��<�a ��j>��B�q3������h@�J��f��)�d��f���-�!D���xv/�b��+���~�q}S���x�g'n�F9g\��3�O}�L<�@�G#���$$K��w�P�6��2I�ޕd")�W��Ғ|�!0Bmx����DC��%95��X +��,J�[�t�/5͜���?*@'���m_)�M���O��1�Wm�/������c�+��0�,�d8�ŭ�ׁ����~(��m',5�=,fRh@4kG��.�N��A�M�c)p�(�B���&�{��Wi��@m،F�|�����*WqBl���=��@_���[nH캺����]p&����19Px:�5�^)Qlo��%� E��7}�4�� �B�SӅ7��`$�����|����w¬�M\~G.���ړٞx�_0���PLY#<�̦����p��} ����ܕ׾�lM+y��Vb,F��ڃ��}��2���J�	lr^���Yaߦ"Ţ�`sFD�Sv]Vܾ&�����_2g���-�A�tuJɣ��L�R���n_ֱ�	-0B๏��>�ɋYq="�+��qb!�X.�O M6���@�9M!�2���[��!Ex1���f�m&�2[��F���D�>���L.���«����n�oS2��Ǎ�e��[��p՟���W8��W��C��9z2�������l�cE�a�A~f�A�\����eU��3��7�QI�J����|�~�Pv�fPq���M��̂EI�p>���޳�4;�������?�c�GC��"�G$�]�%ڸ�"����ԞOu6s��n̨1����i��4[�9�2wOw�U�@��l�� ��c"��ي�y��U�P���Y�:��4!.�r��������B��A7�y��?>�$��0��s���;R�K��LS��GcG69a���Q�JF��nD�%i����qwǔ�kJs���������?֩��_��Vp��6[1�v��ԭ�K����n�@$ ��h�Bݘ[�G ��
�a������ԅG�ܿ�����HǶ}��ȝGS�j�&�� )6yej����*�=�����������WW)�<р�e�1��6
�rfJ����4�eU�P�*��0LZx�][u���h��͕�j�4ܪfZOE�o~�$3g�S��I^n�ݬ�f��N��K+.)��C!��5B\x7.���;��f�2���Pp���x|zڀN՞`�풂�J��H���!����X'g���[5ʾ{�U{�����Q�)��k�
��ɢ�2b)��F{S"ѭR�&U!�*8��7�J	����o*:��5�]�2�vL&Fx%թ���Z��l?�o+X�u��Du���4���Z�o�V���$�Z�"��67�1\�(	+l��9uC�B��UepÙ�Ya>��">�nZ�m㧾�إ�₨ڀ8:x�Ȩ���%8Tz�-����8����+T����LYW�ț~�q`[v����ܤ2��E��c]��R}䜅=��挦�͈����~%��l:
���e�S�t��mR~J�Ĩ�e�9�P������[�Fv��^\|L|�钦[p&r��
\��E~Ls��}�\�}a�S\/�f������ 	�oV�O�m]�(��Or!j=�ȝ�8���9Y_ܳxq	��b� MEq�t���~H��������	8���Ŏ��2����j�FOO�(Sm��Z3���p�f�{�؎˪�^hʬ&o�D��{	�����
�t��Bfo�YK��vv�mWm��S*�ݶ��2&�wG��[���]F�9��!�}�Z��Fb��QAr��Yy��y�ke�O� �k��J:�=/%v�F��}�A_��?�R�R���!�y�vTKH5�f�k����|��p�oN�����@�B�/Rz�s	��)��#�W��x5�� Y�s��U->�q�G��'}���k,_Gm�,5�D!C����GZ �$�5��|��Cϗk�dS��B9�(1���N0�˕�
���x��h�
���Zo��.�.b]�v0��ڢ�v�~�V���Һ6�=�>A�q�F����(M�c�	��h��;�������d�,c2�O1N���^����tt�߹�;pW$|��d+���y�2�P����)4��6�����W�����?ϝ�G�N���I��� .�r,$���$���V��F��X�wY�uMӚZ�CF�R�O$�R�H�m,FOd�r�Oiw�CEN>m�i���0��(=ۇ6a����,����h��4���zc}6���v�#0���׫ӖA5�� }e���N�֦"�;C�hqb[N�.|U=��&���n�e��O��=��e|0�Gy�����z�
��n������h޾���!�. %5�b!e���	ou�ʆ%y<9y_{a:Y�x��� �����s@8���R����S:d����:/%.�2�r�� /��ʥk�)1���o+u�,����͏�<���`�a���w,��'ɱ{�[�-k�8S�[�ک���{1�����Ȓ��Cj
�W1Β�aچK6&}tU��i)�>Lo1��zjjfB�b�	���{�W�� )S�W����\ʜH,}�uTﶰ�T��3��$�a�J��-b��3O��E�������BFvW��%�2gZ���/HF�������=�Y۵*33$�)e1����QtC�+
!r]٘f�r�Z�9�	��n/)'��Ýj�m���a��� Y���{ȋ�c�����!��PW����������wi�>��e�.[)'��L��Ӕ�@�ђ�#�F~KQ�=��r�3^���n�XO>�k(���[3����d7ڂ6����ڏ$��%Mz�B�p��Q/�����#o�T�
{�a�A��f+\��!���'��|#�dV�G{� ���UQM��	�T��ʵރ�=?��Mz�h�����4�7�X��)Y8{�m�#�t��܃��k�.�(�����*�#�5�gH� ����hk��� �*m�������l(��y8H[n0HwNd���zZԇht�U�7�0�*7v�����N?��H�ԫp��7����'1$N���K�468w�%?�0b��z��@U*�(cY�q��ǌ��R}w��=���9ǖ4�}4��S2<j�d�~7 H� ;�����D-��}�}pwQ��i>bɊG������iJ�NL@a�F��0Xr-��0�?� s[�<C	�fND��b<�;��M��LS1)�;�|�+~��{7˧�?BÎ�r�ϥ������D�2A�"~�V�r�~*U�,���4��5D_�Z!J��VxL_HnAU� Mg�:�B�f�y�=�o¡����8ʧU�j�:���pf)y���(X��dD2b����{&'9�R�*�T"���߽)�_�w�mۆlB�q9mV��ֿ��Md4����i�Qy��O k�ic2L	�KT�����ɤ��'?)�Je��u%B1t9<����Y��B.�T[,�3�r��Q��F�� �u��B|��:���VL��)9WD
��O!'�g��b��e�f��*�w[Om·��Ƒ�@5��~gt�F��7���X�����5�c%�������)�e��j m#���EI՜��^�m!v���\!^U��W��~X�18+_4�Ӓ���<��f'����2����v���~�'�(<ptpa��)��4K4N����P��=p:}���	CK���eǂ��`������������Kc
�d�F���n0}H�pL<J�톼 �,��q����պ)��Z/+���,�/�#&l�v��.�����[y��G6�!x4�H�K�/0�o7��#�:$Y�8t�ΒW7��/'�^F۟C���RL� �yɌ��PM3"�]��Gk�Q���Q�:?���t�1� mDԿ�)u\��%�:��t��@���3���x
�rzq���4�$M�??���ÎҦ�:�Nj�����z��Z�����[����J��5�x���y�1����A����A��V:	RP�l*$.�X16����#�&�} ����z�岘��`~X6�jp����2����)s(� �^��ug�2�<��uC�����g��τa��%v%�5T�ۊv�@�h��Q��$!~S���������^�Ƅߢ���T���21���:����|����=�~�c1����j�.�e�J��2�����đ��P��&���+^o9XdDv�����tړ��t�Ƀ�X���(8?�o��L������۱�t����1�Y��:~�!`��"�r�0v���mv5UJ��s˷���.�2��K�̯|�QI�لb ���(N�����MX���ڂ (ju����S��Xl�,���L�_�<��n��"Oj��!���Lv��k����r�ǅ�����)����a�x���R�{�]����;JE�7�$TeD2a�
�������y�]0�v�t��QG��H���;�h�X J'�0Ђ3jLs�s`�����AvL��J\:6�+�^����w�#q�s��� �%TiI�\���rű
�j�T�
�c�5Q��nTe�t�W����9��[`����Ab�C�3Р�Yԕ��s��Q�1Kg�r�R�2~]ts���o5C������3�ԉ$m}��yA��o���?���K�M�� �݄�>����ڡ�"���3��h����{�#�\w@[��I�AߺDv�����Gѵp�"��k*Oh��=�K��P�&�{���f]GҌ�v�+!�樐��ChR/�Y�Q%0�J�L۞�����W���Ѳ��AQ5�b_*	VT�-���b}7]0��$�1��1h�,J����i )P��V�O���/�� ֊�%�0�b�ǧ� �wZh9��e.=p�6�y�a�2m7�Fޠ3YX��!.LJ��"2/��%_���(-z���%��<wF��JT� �W+d4-�Y]�M��
�Q��P�Ө��,�,-I�
���<e�px�Y��y]4VF1^\�Q�ڝϿ������*��F�^e}l�����%	��'(�XRT7�$�b�w��g���"��ѽ�8qif����l<.�H���H�Hbk�����*����L��rF��b#s�u�3��9����x^N饨�e��5_�C�t后{V�m���d
ty�F��KF�U��saꪨ�Sc��qVAf��+,潽a�T��%,-�f�� /3D<\K��~'�9�/f�E�neM������ �]�X��f5�O; �U��{ͮKmL�nI[�/f�A���}h��ޅ7XH2OlSɝ��1�7��5}�WDj{�^`+].�;���1S����w��@9@x���t�8�q������H���70ug%��T+g�hI1���r���L��dE-�[�0�[|I`�c�b!�<��J��54��x�d��&20Yayq,�']Y^?����DB�yѵ6H�
�R��Uv��]�	�	 �u��c�R��~}Y߽�ۛ�JGk�	L���ʵ�/�¨�;�J˿��_����\�x���=y���cN��_Y�q������oP�5�ʊgOa��e~5w��J�󟴈\@�Qx�������S94Q�X���6'�q�Qos�?:��*�	�iH* ��H��w r6�9����p������4��:^(��d����������R���m�6�f���`����{C�c6W���f��5��h��)��A���7W;���&����&��D/�����T��Z����>�_+���/�R����.%�Yֽc���߯v�j..K�yU%s|����lb5��*��}��U�#Ɯ�.8�G��g�C{-8��t ^ ?�K罖�C3� �g������l��@5N���"���F���f�I�rw���,�}��}[X��<�)41
	2�(��~�3��M@-�l���LQ�2_�d���L8 �mӝz�<����7��h�f�#�D8_8�����r�@�T��R��U=;�����8K�&����|�nfh�Fuc��N�Ø�ۅ�U����?��N�FiE�H��'��+���h�J��3 -�ٯ���a��'?XN!�}H<��/-
:!���v�86~\�r=ҠB����`�K�E�U��7�6B�vH�CN��:Vt�;��4ԳU���i�r�)��~��������R
��`v����p���i~ö�48%JP��.�-�)���7��˒U����,� 6~�v
u��'�
ï"�����Dai���^�|� ��(P&�3W�]Ou��?"�o4E���qqE�??���c�ۛ�ʫ����¢=�q�T�E[`���Y3`��ȸ�욙*�ݨR���M��Q�c&�����F`E�a�E����o(�Z����7�b}�;����&����Fe�x�6b�`GrK�+#Q�Utc� Bm�x��*�bm� wA��ik��&r���ѧڭ��O^
��;�o]>�[Q/ʎȖ|#_���Zڌ�ϥ�nqd&�o�)�a/��=���	��Ǜ�j/�A��	�����ߠ������
Tdd�w��o� �)�o���P7�����R��n��to�eg����{��G�v��R<y%���4tA/v{��UK@J;#�k]�������CGfN���$�n�ǆ�9;VVO�;��~_խs��XZ��I��h��1ʈ)7yQ��,N��r�
ۖ9����<f|M
�2�WO(@Oac����9���c����WLm�l��{�p������E���4�d�yj��Xޣ��2x(��]�*%�Y���`���!��f���s�����}ܸZ�ħ���\�m�˞F'kU��S��ӟe }0{���[o:�����uUy��kbw`POm2���������2<��(�Q�6�����r�4��^*vGVy��,��%�d�	�H������ü�j �2��*������}}<��*{��^*zķ�)���ۂ��@����Ň�ǯ�Y�\�^D�, ]o���n���#(Bؗjm��d_W���5��T��w^�-Sҋ%����BJ��!p�D�8h�B��k���=^���m3�RN��T9���?�2����H�㿌��6��R5�O�Ҋc�M @�<�풲DZ�_l�x��S]��}�~��<�ݖ�aܧ��A���Ԓ��έp0��d�"k����?F��,���"g�s��@�䐀I=1�6&�q���S����?9�1����}�#�S���h�+���ݑt�PH[)A^��.g0a��&4r�s���.,'�zb�*������ ���<*R��%�^}m]}II��'x�Nt&E�9E#!e@Df���;�[�b��d6��kk/�Ѐś��/�|G��f��m��}4]IM܈�U���x_U��pg+G��p�����U�"���H��Qɨ�آ���I�ݛ�j�*^��^Z�Vh����IIl��p�E�%����5���._7��	Z���2;r��t��a
s(8N�/`�t��W|�Z[���	�͝���myp�=��
������<B�������?�W�ך]5�&x}7R#H�st�S.��w��9�B˘��u<��nB*И��^� ��~�zn�P�/�CQ�����?�5���]զ�����m���n�����d����p�5���F�� Y��w�n%��Q����6+m�����D\��HGhU�ͯMKC�]$`!�� ��3�A�Z[v4,�[���;�w���il����Nn���n�>��6d]��Oz6�3K<�0H�k�"�3���#���J+L�&�mx����h ���g䫆�a�z-X�����B_�Q�L:h W����T� k���8<&68w�h�K�nhD�_lD�<������A~8��orh�@��y�[��T���A�x7
(H��=BF߸��]6$IՂ�����C�DR�,��az���}�^.y�#�k����{�ث�U�~IM���#�'(��D�H�5�����#��7�-K^���^�����\�i���
"��'n��rVF����f�Q�6���/y��0�#gM1gV��"΄��Zf���aT�-�n�����M�Ę�b���jwر��]��-�����ޢg�+�I�mn�{`Gf�[5�-�s��^�!��7N�}����|0%e���/�V�F5��o��e&����Li;�B�Ù�6g{���y�����_A����\�f�[�!�&���� ��؞$N�	`".��a��S
��G�粒�HҠ)�ȗ�p��hW�F[~�2�p�Vr}�0�����-��a��:wk6�_*���'}�t�s(Eg��A��,��ɥ�x��@ћ`Hx��44Ibb^O��S�57VP�2R�`�KFR�r�cK�aNf�ǂ��3��V��V�҄��K�#od�c�
�&���4?�ډ��q�һ?1%j�����]&�����{��г���v�y�U��%�� ��p�#����Ml�0�����<��)ٓsNU0a:*N�L����
�kY7i��T��zँ�:�4ҡk	��>N<+T��y%1�U�M9�e���yZG���J�u�֊���2���Z"�v������@߯�I��A����ޒ�ZR�����Ċ)�聜`�w����h��w�FY��+A�27pe�?���������W�m���{ �5��4˙�����&W����Re���~v��Fs�Tf����&�ď����� "����e4qB��b�,�[sX5�th��K$�#B���j��@o�]i�-m �h !�g�e�@��:` $j�6��9y}�ա��1wA��L����ر.dn������)`I����b��������C����q���2�l)W�.�*�rz朻b�]�3w�㮳��d��'
L�m]�G��%=Ǖj� a���4���q6�C��c�%�}O�Y30���X�4���h�Q擄��)#���Dz�Sz!Y_�b��;!���Х�h���4�W�6=;��]d�-{�%ƇF�G�����P8����=��ߦ��]ŝ�[�;!��Ys$�p�`vϘ Zt[�TVa�@��AI��p�\����'�1X�BZx����	��wV��v��,i�0D�ņ֒|0�fr��}�������Y�>$/��pI���6���Ҙ3�D2�%�|w�4��4���mX����nhw�T�Z%���f��ïV��c�L瀖���Bԡ� 9#�*����O�Cʴ�e�Ep�x@|-PN�"��s�9ע��2�ƪ>�3�"d�Y��1�I��{D�rz�t�$`�:�ڂR��2�@g��\�� ��v�ɋ����|`��[�w�\s�}-��5ȻK{�?G�Z��<�D��^��I�E L�
5G�B/ϑ�!���=@��LJq�ltۖ���#�5��oMF�4jv���¥{i�Á���6�e@U����{2�rg�~�uN�V���ck�eN��#������F�+�\�#{��Yr>��B����H$��+�R�>x���q�F��,=�s�L��ORqn�!���	��"�;�5�:a�T��F'NS���� �n���5��]w�� �4F3W���?�X�y�A�׻����F||�D�;GCP��"^K
��׎�0ȕw����rE;�~?#L#��u�7V�����t=���G����;���&	��
k��OɌH7�F{��>�.TZӂ��a�ܠv��d�{����,-*
���?\E�E�g��)���:NT	�д:�b����.׹3�̠�xX��2�}!0��@>��J1��[Y���K�Uc\��n�+��M�,�F��V�)O�R`���Q��������A��(ۤs�R���$��d�K����2JK1y�%�B��),�:H)SB+L]�Hc�'��IKjrɮ[�I=�V2�]{��K��I�Rq��m�^�=_�BG���鉨�x��$�n\�a��mp��G<I%��$�h��#P���S�s���&4�z����&e`��U+_r�ݜB��f�5�p�3b}�`*�Nk�%�{��+H���(}�1��C96�-	��
�l.�sa.,�
N�q��3����,⡦��*�p֮�C�*��`1��t��u�	qjĐ(��Y6[Y'�ٞ��� "�w��A��,�{b4�մ<��M۰ʼ\|��P״�a�e>2�f� ���H�\��|fzrfՋ�C	0��D
� ��0F� �f��>XQ1���B��p�l�"��P��0i�S��
�j[(�e��+�Lg�������l�A��w`$���.P�Ց��u&��\Tk�$�|FmLik������� �gX��k��[��b�~�(X��ī���F��"g,N[��w��Lww8�����M`,���hG+U�BmX��AЄai>A��!���2'�ȫ-�^�aV��j�9M�'
J�Л5�s��t�J9܄s\ ��j���IE��-c��X���FI�����z2��n!�9�ۚ���wm_+�)�k-��EgAS���h���9�� �aQ����s:>��-x߁����](�~7�H���y��:���#�|��l�z_B�\ׅ3�i�3��R�a\�4T\U��g��,[R[T_����T�);�J��1�҅W�gI|NYo�����'qx��nu51wʟ=�'�~�V�[r`k�M��{�/纤��Gt�IM����ه2B�p�qN`o�{w���e�7A��!��Aࠤl�^&��wP��E���e G�7�y��ǂ��-�g���{!S�
�<*ҽo��(��[��$X�;j�ʐ�iv���̐v�m<)�t -�
@�r[�4\ ,F���{�?�8� �O�s#J2�-i��!a��K8���^��i+Vӛ�N�t�X�`�HaʖƧO��Q[�"z�i�AN��g�* ����S��8�3- �1-�Oڥ��\pk�4,r[Q��v{BK��i�Q�:���� N`��l���İ�e���Ar��#�-���T��n�K�9�:bढ़(����s��Â�m��/�E�&�$5o� �˫L!���l/�4���B���ȝ��)3t��H��X��m���_��A+!w'��#�:�*g��^��<��5��CkCr�d��lm���n��w/p虧:C]J��>�x��(uw����S��G
74zl#�S�ErA����qH�E�$�[&�>jʔ��Տ1�P9�9~7P^g�GD�
��X���x�24��In�OrA�8ԸN8ڲHH?���ú�6���Q]�
D>��Hq	�#x{JH�k~W��*�n�6>b��'?��CG!�J	�_�������q9�M�T�Aig^7��� ��>�Y������.�>�k3�������0ߵN)0�^9�{��w�.�m�j%T�d�Sk���+|�����ϟw�7����F��شo�%�٤���R�� oMe���@{���98ݓ�Q`��`���IQ��j�r �}�,AM�o����f3���D*é[碣=��p�q�P��^H[|b��	�^X��Ƒ&<��<7=�9|`Y��I�t��؎R{�m�6�F.�.B#�TK�_'h��W����B���Yb����.��y�<�
V�9��Ɏ���N��`j#mh�V�V�����:�F���z��<��Q��('�.��t��4���#��&I�Tz5�!����������bt��;�����epK��V��^���Ǳ#^6�z��	v��0 ���+<$�b����M�b#�s�S=~6�W:���y.���qL&��I��X< ����rF"��Āa�΂�_q�����23��<>�����ж�s��dm^\z	�H�Ѿ���K0���An� ���Θ�HS�� 1�dÚR�=�墺P���Z.$&�T7�V�YTɃ��;2f�qo����u�e�Dw��0f輢��h�BG�`񈯦�����+4��x-UҪ�P̅6��Y��*�<b�|�� =����� _\u���U���ߪ.Y�P��V�U�L��h�|�$ o��p��*�M�c	�S�X�F��-I�ad]����Uk[�K���oT�����쭋`�*h���o�	a�sS���,��%� 	�6j���5�,<����P�'�17�By8���5'�3����O.</X�Nyw��T�/ڪ���l�_�bz|�gW���*�ݏN��x���p�Kb'd���X;x6ՀG-�N0(���N�c�`��%Q\a~��i�-jo��'�U��z�W�Ѐ)�1t�Ns`��� &�ɱ,��k�����b�������+r�,tn����L��i�M)�;�:z�]�J��k��0Ħ����L#B숟��syq�*�������x��]�&�9�g��<��M���_����w�5$5�[��6P}�N�QЫ�ˬ)Y˄�o.7Cu9	ΚՂ���I�L�i~�g([�.���mL\�l�-z�����: �-�~�+(����2��'�"�K��T ��=��-�I��@�q�ʼy&���u�#��q̣�dַR�+��X|��꼎)��قܳj�\��NA��nd��<l�.��� V(A±��ұ��8���O��C�`����B�M}L.�U�Q0P�*	��N�$#����us���D-�N��V�)��,���"'��C��,��Gp��� ���r�N�	t\=�Ŀֽ@��ďD�^=��k�pp�B�(�o_��S	L�Du�S9��͉�)��_�[e7�<��y���p��s�Q������1.����g``'F��Y���D�3(�Cs���5@7���e��Dv�Oy�+	w���\2�Xۊ�k�hn��W}̨��S��l��a�O�`~/a�"9GE��В��kl4���G�K�[���@^!�+[��@�����j`Ʒ�S��!�v�����ﶃT<�n�����I�i��������L�K��
�m��K.�<b��^ے{b��d�h�7��0YT�!Ϫ�I�r9����3忧���ޟ��Y�%�s��ǽ�6��Y��ղu�ɴ���׫y'b��Jh���.��=��#@K�[g��x,�+�=�y���X�c�iG��:�*j���:/I���G���6�$��G*I"
X�����C)D�s}Z�����n�H�Y��
�{s�ݯ�)����q�L)x�X$�"+���������[n�]`����5�y�;�=ޒ�6Lҩ�;udA�q#"�>E�����.N-��B=�㊍�\���0��{yO�3)Ja�b�M~�DӿJ:�^ҕs�fl�*=-�ytj�vH�+�2��jgC_��'�ͨԥ��m�1 Wɱ8Z��y1�"�Ej'^D�l>��B5n�}���OrS��!	�l)�M�Q���&EJ��%@����s���{q��ӳ�Gq�+��iE���ț�BDPV>6�EDT/�FF�P-(|����Vw`h��2���{)��BOrmq���D�7�(S��Ղ��P��t�_�P��t�Pz]�"'P�ؒ�e�`�'S5��12�gU���=ǋ������l�Ȣ\Po�x��hgO�&��{�����,�AAwgd�bdחvO�H=�'���n�q�T9Y.|3���� �~�aP�����D�(Kᦍ�5�S�=�H��{d\�|����o��w�T�/NO/f�7�#$4L-�;�Dd�!���@�����wЯ}j������D_(yR'Z.�rg@;\`�F�bٿ��}aOBC����N4k5��Hm����	��(&k5=6$FB�ⰳ��>0�hg��J��Z�ciҸ�ߟ���O�T���?kr;SZP�4�̓���"���Lu��5�8ߔg��~^������@�&x��4LDO�P5�zl��XZ�țZ��/,�;_�GH/�[��#:�k�~1١��V�C3fY��fR	2�Z�f�H&��28����O��Z)�����K`$��k�HJr-$n����û�X$�J���'�8w���U��e��ȑ<P�nC�]����>�@z�=5��Y9r����T���0�~�2q��������g��3�u�Y����t�U�����[_CC&|Qz�U���Q�%��������#s�n�����M�?�&}�-� �#�C" C�
23���5���A�`��?=@Ye��,_�B^��r� DQv� C2h6E"�V�z.ޞ��m!t���޷���dm�-�����)'>5VQ:\*uCqt�53'�/g����2��þ��X2�,��zb_]7��Ge��f ���O��f�#�}�tK"���x�IX�8O�����q&5)0�~5kP#n�j���#"��M�&F���YP�R=���#�G���r�~=�+:�v�W	�Ӑ���Z#�q^�V�[��(%0�n���~�
F[�� ������[��0���$����)�^�����B�m��	]�]��>��;��t�	k�.u��x�_�1引��&U�_?;1pgJ{X*�S���w	Sa�]�l����C���8*X��U��U���:r�A�U;�z�6�.��Z��sC�3pNr��C|Rs�t�,��F�r�ԡ۱����`c5Ha��=��v F���K(
U�����}P�L�a~~PJ	9��*S��uqct�N�b���g���D$P o��B��M-�]��s�����6>j�>�"ۺo�Ab�ё����.�~J��
��M�,|����
-�ϵrz`i�"}��((7�N�=�\U	�Z���.^�;�1i������6~��.�q7'%�gΉA�v_<�Vg��<7YZ�}Z!��ēr�k��צ�^N�
�ʥ��)����	��������?TrG��.�;X�'�i_�%3Gb��c'j��>�$���(��1}���<�:R�Z$�Le�eLF!��Y{�+!lߔ��{��s���G�@:��⑲ح�Rp��n�8Cf`���$ӊP6�"�x���'<��>�~9�� �=�l��j|�pᓇ|��O�����)9)�E_�"a��A���B�S�IB?���ki�2jyB��#)Z��̰t}��nP��%��Z���d��cqJ�/uh�����5�t�,/�������81L�z=p
 ��!���� T���U�Ȼq�.�;L&��FΛ�Zn�
��DdK�њ±��H,cQ����_�8	ryJ�������X��y�Kw�z\�[�"=�EI�bl���ԅaj �K[���옋o.p�͋�?�c�#������ԉF����}MzG�H������ib�	���p��s٪N2���:(��漖�b4����;�]Ѝ����<�`��)�����،q���8!��ٰ�#R���]�I��P�#��:X��� h?c�t��$Y�<�BVݭD�J��r��4@�j� >��9S)o�BU���6}�H<|�B�SA���DS& Xf?�!�ː�+Ү�k�B�������05���Y��n��Հ?������4����|�J�_�o3{Bs8��#�S����[SA1|��b�������T���^`"̓$���S(l�t&L���9.$�0&�d���==l��ҁ�t�Py꠯ �z��#^��e��j9��h�K�A�`J��{���A2+�L���(׃��H)W� �2����@��Q���톣Q�����i�!��X0�ʒv�?Ț������Q+��\�|B�d�	�#S+�jfh@�P,g���L�M��fs����TP�A��tl�idAB����M�E��I�D��R�վ��}s���0� �|d�`
�5��]��V���@�`��b�����f����j�.9�\��Mc���b�^h*�l�a�.�	�O�qL�ܥa�t�j��9��np�D���Nd��ɧ@laƁt��-	��qȼ(�������4��"x{U�Ñ�b�a��qr�È�4��^�c��J 5���t���/��?�ۗ�O�P��GG6y�x�\\��v�Q�n5��P�Q5�zI�ㆽ'�����C�v5���|�0�*�Ӊ�Y�[;jA���P�%�K�Э쾌{���G��\�Y���V�O��w�UJ
O�4V_��+��6Ky7$ֱ��Q�C�S�*Z�j��;�I+��=�Ɲ�Y:�TG����/���M�y��^_����;M:��4���N�9L���w���\!���>���g>%����úp9Ӓ���9tP+���*�Yj��.�}��s�oԉ)�����GR��@���6��/�9�?鰧��eG)|�fx!��X�(b��	y����8�A���5�TMl�kH>ړv�k�xPt�jHw�Iα�p��T��՛0��o��|�s[���Uv\�V�L�ؙ�Bm���:�z�Ճ�$�K����h�2�C�4��ņ`�^��z�")G6Kꇘ�{e�c�p�M"�rF��o|��"��}��K�!8��v���lQۂ��-�M�v!���*�4ؗz�t0`^�@--��x۔���:ʢ?d�#�t������#�Cسj���)aDW�>ݿ�&]U�5�^����B�6(>`Hݘ|�/�38�ߒ�d�.E�� KV"��v�W	|SZ����]0�&D�d��E�Jh�l4������_��+��Q�qTDJ��۹���k���4��"q3��AN�uU� m��^
eՔ ��p�*�ŷ�NͥãWSW�[z?�ׁ��ף��0t~[�G�[2#ˡ�̥�_��(��p_>��~�Q�^L�f�X��!�	kp6O1w����\����g[�c���m4�����ޒ�p:��asb'x�.8�ŻRY�X���\�u�u����%�;�{t� ڣ�m��*[�rG[)0fY��`Y��\���_B�{������
���L↓Z��̓���0���e��mM�<��Ĳڙ|~
Y9��,rp=��.5S�U���ǅ����^�?jN�j�V��t�
ˉοp��j�.,��l�p�U�M�껰�@z�Ѣ��j�KLUtn�Whb���Z��U�9��"'1��;�.��!�����+f���p�D��!w�.yt1��Yg5i{���N�2�3&ÍY.�W6������n����Ϛ�� k�&�N�������b�t�� � �l��m�؎_�{� lA���ɉ�:�4m�f��Z�p�$wU,r���!�(�! ��h֜*�x�H�#���s�I� g�CX�����'� v�Je��x�S�/�0�Bۛ8U�HA��Y-X�Z�2pe�#��=�
d8�5EjzK���t�a���"���FD���ǟi��ؓ�z��G�|��b���������$��B�p����p�G2�.:���O-&N%�b��u�Q�qA(3��R���I�>a�C���6Rz5�Q�y���;}�cyL��ѭ�b� ?�2�_�P�bMD|݃G�Z�ˌ�B`�tx]oy���,]r��V��k���e������6����?"?��	ʻ��v�ة�{��6X�jg/��o3�+٤�^�~14X��0vq��� b9�7GSc1�k7k�����2����ufo���-��C��$:5�=z'n��#��18�&E�1�L�:��ĭ��]�п�m���T	����?�g��1��(���U
¿�C���hg��>����9/h�e"_O��P0���>+�??c,�B�*�t���=�>�����dF��zb�s��3�$т��rȃ-��`�ܤ�K��:���`� 3���!É���8���KU����0\zi|B��p�X�u�����҉x��;�2>��{k�´���j��A?Q�]����{��}y�(��<��IX Ǻ4���s<��.���9ܒSܹ���>)�C^��*q}��+��>#a3��1�1D���) �rh��LGD8���?7��[�*��>�r����#o#{b���E�F�V	��6T^f��Hmz$c~�d��~}�K"����1��H��_�{y�KW/w�oG���ɢn\�/�3��ō��g)��(�"�$ۊ�?%�JEx���?E@?A�w� 
�R��C�(�K��jR\�`��}�G���,W�o��|�!a���S�rӻ��nM5�M^8��|k�Sq6ȯ)
u����P�������$=K$;��+tsbEac��;���ï�A��DD�j��G2�@X�m���cNn�-��cW���WPʣ�J�l�j�E_��0��Z��*°�����"B�V�������m�0-rNȈ������M:��5 =��ne�S�?3�A�'���g����v�O<�;6�%���V-�*��TQ����p����Hm�N1�r�Y���W�tSGz��!2p� D7��!{��?/){��H4�T#���׸T�Z���V1&%�"��H�"Mͼ�߂c:���&58�ߒ+ m�u����u� �AW�,�JǨ7;;���JaN�f��v���g�P�E����~8�)i���/�P����"����Z�T��ں��DD�?��l�����UL����M��Y�(�F[�w&������e�FX����|�r�G��b3�V>=�bu�m5��H^��=V˾��.Y
��~������f"V�8Z��n��d}� �d��~�����t�{37 �3�Y@M!��M�����ֽf�D" å�	��O����pq�Ck{���
cl@�o����Lwh���,��6&���+h�ŏ����:��Cy�(�LF���&�m�[j�K&���|����K�麅����5�(Sz��Y����ۉ/��#p~�^�7���i���)Dl5���3�6��
���YL�)��%��q�j��j;�?r�Dt���G�C��$<?���I�����?�bRF@T�#�������A͟tq��E�rX��A�r���`�$��1��>����n���k-�?N?���:?l�%v�B����EL�� �7;H� /�P��)W!��24�г�i0Ӷh���&��`z;r���5c�Mfߚ}�`��N��o�7g&�I�%�H1�yXcJ�_���+�����bT�D�Բ7�oi���/�j����R�2�Lr@n��!�lo�}�835��|��F��<o���B�C^�3�\Ϲ�^"�l�B�D�a�q�rw����H�sE&�����@�Rh�-&�7=,����d�[���^n���[��_Xܜ�	�.%"��j{��[J�:M��o\��}X��:��$S7��FEKaЕ�#ɞ�j�P���94��o��OҵY�GǦ@�[YiSԦ?E��~q8CN��L�\h?m��rc��
]l��|!@�G*�����GIk��Á���΋l��5�F&��@0��I�ԷL˔gc�~�����"^(��զ˦��,���G���ѹp̖���6�=Z���X�ݛ�X�P�����n��b����!Z�բg���C!K�֑<S[T�7�k�ײ�����*��~vs��_A���90�y�+�r|��R;����T	�J�"SPKI� ^�Mnf��X�%m ���r>�{�W�����8�򾣉6�̞Io���I�M�b0�|��^�g~�ک��yB7N��o���ہ��F+�T�Ri^��K`LS�}~�D��P�*[���#K�y��4�M�P��r6�2�o�07�E(3Wרq�y�}��1%���� ܟ��h��Sub���vѻ�w����p��wiDƍ}���Wd��(Ґ��_���NZ�
�J'Y]�W2i(�|�cn�?K��^K�=����{���pDa/N����9����@��e
�>(��<Q��?�!?�)o��՝�����-�_s�Ѻ)C��:L�N�D�<<U~`�i���}���g�wO�c:��CE�B�=5���5�T�eP�Ω)W֔%B��0��~��}X�� �w���۞�B=4o�� �3�H?��H���)0*�/�dNW�Y]3;��<�����X}��Enjm� OJ�������~< ����:��@`� *ف5�i>�+��h ���k^T�8�|���oĳ..J�_���"k�Y�`}���g�RJ?c�1�4D�T`�΂/���6�?���C=Ce��`�
4���]G��D�uy.�
�̘[�ET��sL�����D�UWִT��[��E�U&m�wu�
}��(c��&s����b�"
����rU%�;�8>�S��h1����~yk���;�c�����c��ʔbt�x䎃M�y_a�{���G8r��_�CI�U�=���8L<��<��Q�VԒqh�x���?�e!�d�K	�Ug�\x��D1B���Z[��7���<��i��"��jP��e(���x~�x׶&UN���<��_�z����ԅ�I�Wj�A�F�U�
�1��p�� �g�ͦ�j.y�Ŀ^�M��8�&��=��rn�Q���|+�i�D�R�Z���.&8#�PT;������w���#�#����MZ(��i���{��dޏx9jW�s�`|�:�9g����Y�x>��P�o7{�ө l��J|�@-��N�fE(Q@<��<&8�xl�/�-���+�(�-
$�_TY@��鱏��X��%�TC��U� ?�>�Gz��CL,��SG�����6�r���6��������V���k��g.����e|8�`.��x�R��U���*\�X,@��o�<�� ^|A�ƃh"��v�`��%=�)~=���;bf��X2�L?�24����k��UPI���/��2�+�g�sm#��ç��q&�(�,э�O�, ���eg	UՖ(�-��k�5@���I�	 |N��I��6T���̐�����0�F�"��`��Iᚿ�f[��J)��.:O��Uo��*X���:K�Hc�f���+kV�~�	��r�V���U��I��11C
 �!u�B(\>��A?e�W��WuR�� 3�x.�ES%, *|���S[.&���K����t13DP���k����J�k�"I���mT�W���;�9�w	z0�7�>Ɗ"��"}o?>�oՠo0�0��@�>t��b`U�M���QXt��-� 8LИ5�7��-*��\�8~ È��WH��j��0�V�4�緻	jT.�kǅ�,g�YfF-�;6D{���wM+�ћ�ve
1Z���G1�=�T�;��	S#A��9��p���j�B���u�GVR�ļ\bx��!:���7+�
ڟ���p��:wg���r����ȳ2[\����������9���p�s/����i�"��c�qIdTw�j�,d� R��`0U�<�c�%yݢc�������X8��]*�/�+�_r���辜�
ƶ�L���C����L��b�Jjc7ӕ�K�@1�;9< �G|���$|x!��P���J�*�q� K�����X��k{`�x�טs�4Q�qc�ί��`�W�ڌ~|)>����O���@��+˚�&<Ϣ#�	�2K���&|N�)�y��:���mщ�hi�6̍q��^t�	&�
�;�4J��3�aG�.�y�p��Xw���_���x����R��d�d�� �V���'VH9e��X	@����C	o�*!�nmK���y�W��K��<y�!�l1?�L@+�wd~�%���|��u7��"�m�C�p����H�S<j�d�.V�wS0;K*)p�)���Nɇ��D����=�f��4�up�eֆ�{�l��?�6��D�E\�X1|M��Ƹ�m;��C�L=Z��u/U����s�z������|ьo!(g����~��<�B|�3�*�PZOp[���a���كȳ����Q���7��;	4�K�>���O0�>T�N��kgn���{�d��?������Q�����(�h�1�ޝg����G�!��G�6}���!� ��1jr����֜_�~'O������@M��Z� �x�dj�4y$:J}ƨ{l:���%;.}_a�|n��fjުT������h|�=6��jT�-���z��24-��� 
��7Gy"��J��(��0��TP)��V4�k��[��@�}��rm�A�ۣ�*Hr�"�_K�v����Q��IOQD�N�~ؾ,oCҺ���g=�I��jrD�{��6�w���&�T��A�z��Lq���EZ�o<'+kc5aY0�L��F	F�ת4�@����y��CN�`�>s�0�TLUN��*Q�� @6�
VK�EY�ۑ. E߷Tֲ Q+�k5Ŏ��5ڴ�C.3êP�v�I讑�AqQ|�Y����˓����mL�a_��:���[��!�'��w�ЍKr��OV�� ��~��������etx��1�^�����l"�'�	%.���Qo���P˄&(lh���]���?Y��,O3��?O%>��6D_;�A���ĳg�q��Q�ě�:�����a�L"�(��D�.\�o�ZcR���m��w�4��y�Y'cX��J��>��5�r�X���+���ܵ,���`���o,�.�t�1w��	#Lq�u/��p�4攮f�WEW�d�e!~�<����h��+��|�?k��}�2��$����ֺ�n����,��2d�Ӽ�_�V&���"π��ԁ/ո�N[��^!������&���_�,�pj���R���ns�X6a�ㅅ�~"{4u��i �Ydj�E�֮S7�� &/�CZ�V�l�o>�8F���+By|�ާ�%;
�A�F��9%D+�3mF�]���aLӮ
����l*y�^j&�ώ�ta6AF�ɴROm g�zYn��B��b�v�ta)��F���ڧ�ʬL���F�����2ts�'�o���F���:ژ������� O�`B�a�7��2����$�'���0e�\ ڱa�<(�WS�8f����`1&94U�UW��pu���N��_z$V�>��n���s�
)	f�`���+%�"��a��-&p}yIn� �@�&0���V�����{^�(x�E��PĨ -�k$ٿx���ŋ��$~�+VOspi��EY�r�&]_�H���m���Cz|*�,�B��W���ْ�[������N���-�������d��+�rq��B�f��ɓ60�	|E�nO�e�6��c�f?��Ʌ�[Bp�#y��c�L��
j�i��7}��D�l)��K:�Q:����2[��Y��K:I�
���_fY��{Ƽ�C}�I�c���b6#��LNZ�dD�=��S)_d8K���8g��w�yBW�G#�,�t8� 3n٘
�P:s,k�«�*��MC1^x[6◅�8��k��.&��i!i���ִ �����`��*.��{в�.W
#�( ����8�E�}%�#��jSr�3c��MG�H���#��0�	��t^0��r׸��'I/N k�9�;�>�m)��r1)@1��1_�Ђ?2�%8��qe�0�2+�:���-������v!��(ov�mN	�Ͻ�������H2�m<��Y���Y9q�&M/�W8�Ptlh:_��Ŗ/�0 �|~-��-�}�^�ew\���X�`�I�lK���R
"�i,|���b�]ݥż$&U�r�M"q�ա7��Wlf5� �P�&�i[��7�O����i�yD������]������¸2*b�W�o�/[?��{_���D��*(B�hf/��^�4�g;mz�t�]�맥%Xg��T&m8���oU� 	m;*���T^�I�1�MҖu��5Q;��u�mV�@����#��ۢ�ȴć�9�cb����A�AhI������ݢC�S�M<��)����tț��<����4m�o׋����5%�#+,�^"i>����P9��w(6E
�ψȻ��������Uzо�m?�����S��/����@Պ��ڮ��"Ȉ=g�qM��ֿ����'��0�!�	��8�N��07����f3��}�-��
��-JT��a)@4�E˾�Vn�� �OWv����0�:`�a�b�.$(�s��,$N�Q�]u,ƍv�Ď��e��3ڐ
��*Q�,�8�qy�Wx�S�&/*�|�LA#|��9^�����f�:?x�!%�"-�4�\ql��%[|����3Z��
�2��.Zt%Q\j��DD�;�eQ�Lü߽�9_|И�Z3><�<�Uoq��̦2��{4�<������vV����?���-�\��g�����n��L�(��0�o�w���h��,�h��1l�Kk��:~|- <�Ӟ�T����Ų��v�)3�!C��!��nm�|6�e��Ӻ^ MM��ޗ��A_�$!�(F<5\*B_Z��rJ~8�P�%��_|6���kM�+�H�}X���>��1$�޽@�z������\)���"�vK2�b{�+�vf�T���*,�,k�v����:	%�;d�W���N��F�P���>o�ě�^��C\��^�o_ݕٷ��F�Мj�T���{4��-��Y�����oir|ܵ ���clD��L�f/ܭ�?T�!^IR;�[�U1�hl��i�<&��']�������~���Z�������͎�+��>���G�z�O^��si�D��A?�3�pԘ���Z��9!8�`^��S<�$z5�sv�DgF��"Z�r�l�zhX��N�G�bv�S��1�=�E�]92r�o��8�!CTo���$O��;).;K-p�f��_�g&�T��	�:�W�^Pe��q��J��6h�Y���h���;�������jԅV0�ݢ0+� ���Jhh��6�ŮC�"ADڟBH³r������ZLH4�=��0hA�ߊ�_�Q�|b/B�u�ؗ���46bs���i�/��R���4��)r���C|���!���N�㘽���i(�����!&b+p�b3)O: ~m���s��Zj4�~۠�/#��6I��Q�4e�'�E��'�:����%`er�B���;��xN�C���#Tb��)r�����ԢkX���ո�Ę��;�=��AdǙ�v>ڍI>�~�IZ��c�@e!ν`��V\D�7�k/���GT�6\w�0	E0Zc)�H{?(����%F��^��"e�H\^�G1 0��*��u]s����Ƅ8W�l�\\<��w�h=�WW���>��!j|ez<�%m����	�M�Lh]�=��0N]
�%��$�r(Uw[���Ms3�y�1D0� �h������W�D��⥔Yn��'�,I���&���M�
�
MG�Z�7��J��]�/��� 
'��Y���n�3s?On='��r�b�S@&n�F�/p�4*�-�\�^�a�aRF8-4%4h�;�����9:n�T���R����ä�\R/��uK���^���DR��޽�67�/A0�L����=/��vٴ-�qϥ?�W�%�I2a栢�.b`Y:�a���l9� 5,��ن����Ęв��uI�s��h��Y�����7�\�iKy�My,s���m	�W�D)`�P���:0�(�5) ё]B�#��m1�l 9���Feƿ�ˊ�/�!{JO��!ne�GI�PneV˽i}�y����nK���' tm�5�^�XV���A#�c�>���?d���!3�T������^�u=���@�
��C��oWT*sB?��c:��f�[+WlmE�Nb`���֘�a�h��#�:>���lyG��ʮ�"�;8���Q�xHI��+ėuu�Cl��ܙKP�5��i����k�hk�����ᴅe5'�Bo��$��Z��Zl����(�L{<����W_+�h��Z�q5MY������}���n��2�
�d����IFi܀��l�X��Q�M�v�.{�'���/Y'��SF�}w,�5��=���ˆ4�߽��q\|�v��CJ���;�h+zF����M ^�$4BF�4�35����*�Te�G�[ �I�(�q�c?����w+t4
�����0�q%�z�(7y����s>���5�:0�.�3�mz��O�+��	�`�2b�XWm˙�xC�ً~���v� f�󃳜��b�9G���(�x�!'�!�%Z�)it��<GQ/R�$г��� e]3�;3S |I�L߽��_'�羗5{����цqß�_'�ٗ��Kҕ}lݥ!�1�)J�(��:�#Sb���+=H���%:Ŷ��
V�U�UQ��F�Z��K%�MB���-�ր��&4����mG���w��!k�����m���Q� ��;#��b��Fw��k�'�B��p��v�95*^���#�ķ2��zN�>��n	��/��q�����c�8���-O�u:C���.��X8���y�E�}�{f�� �Tp�Re:)�Un6`�UK�J	���/Bp7f���"<
��J �����8t��F%r3h��-/St�C�辡5E�4!{3C�/g�Q���_��G�6X9��Ѯ�Q�2/�v-�o����s���T���)��ʫ6�:������8����.2:��4 G.4�0S�!���䰗��Au��᎚m���UN�~�,f{.�����`S�O�����R��'Blך�G��������6B2�L�4�AI%�~ѹ�.����%�P�
�^�*'�z����L:�3�|�f�&���������(�oXM���Շ|�$�27G�U-g؏�����
MW�N��3��y��!vy	3<�F�SS]&F V@�]��%���Z}�Aो�}ʔ;o� ��Ԕ�-)#{�.l��0�ى|�dfp/��㈏�`�|
�V� �,��MЬ�(`� ����C�$&/Jk�	I-2O)kN�!ZZ�#�k����Lc7:{i$�g1 [�8퍠`�,���eb[qx��e��R=z�H�p!�#��z*6Y�Q@<U�Y7�3���ɝB�h���@\G�P��1����YW�2S�6�%*��7F�Vu�6d���i6��Yܢ�h��-p���"8���F�P����Qz����E�XM[yN�T@�;2ms�t=F$�9KZU�	I-M[��>.q�Y�زhm� q�}_7��<T!��������^{Q٤�cg�X����xWspR�b�:����o���]�EzM*�Cю�֘�G��n�<-]����Q�?��c �(��O�j�����Ĺh;�;���
R���A���P6`�d��0���=�Z$ՏZj�4�٤��;���N�.�̐����!��0}�W�Ĵk�q2�y�z�_87�`�#��?;"}�YI���JJ_���LMK�M3���O Fpe�����vE��o���n,$��л�i�1C�9�!�㉴�mHd�Gy��W�DRk�.0L��:Q�Wg��ˊo����J�`S5���2c0�t�/�5r���$�X�;�����
s���Se�)���s�콲��>O3��KTa�Z�t����(��2--+���t��b����5����	Ipl\��dI��|!)���������4��r�O.��'��4����䛩��L�]��2@{�|���E@��ө8Tx�D���f�n��3?�@����Bp��SM����9��6�s�a�����7��p�����$n�8*?E���ݮk �ꘌ��m:���7Va��=�'��(D0	!NiN�����Eܘ%b�O������<CAQ16���Ld ߶w���v7��n�+�g-�%6�~%S4s���yt�M�Ձ"�t��˵��0x���R���i|��R������7���
[e4C_�4Q�w��5�H�ujjz�Mڟ�ʿ�)��F�wI�pc�F��A�scЉ�����Dm&�/A�⤔��Q&�H�u@PQ	�έ��'�^��l�4Q�P{\���.�Q�����-0���X�~$�f�h ���]f�P��u�V�]
˽gte����;�v	u�J�R��<#Z���Q{�j�9��h3�nA�
*~5fe�?����~#���ڇ�A�M�&k�[H�6��y��Oy�C��Q��"s���f$�7��o�S�N��oY�{�~x��;�&8�
�C��)���9�+�Sюo��"��r���)ImjҰ���� J�)YiF.��ӬQ�>2�Mʲ��pD�H����D?@�yB���xliz]�$)S�	�%���Y+��M.��`�\�A����OS kK�9�f]H��Wb�Bf���:VIZ,d�cF��)���9Ү���2nۧژiv"����`�Q��[�A��CA��-Y�л���Y`�^@P����@$3��e�-���'cl�����/�M��� F/󳏪��`Nj� �v؅�<~-�\����5�y�f0@jN��v��Nx�� 0��>+r��sy��{Ļ;Hߥ���D]�<G+�'��\n�P�~�n� af�
'�]1ߟ���u =���cVY����8I�u�l(�ҠarJ�>���`�y�+�/x=��Rd�jP�]4�z��X���L�E=#�.�W)�׬� :�|�kk,�[4�/����Z|m��E����Y�c�,�F4�VI��u+�@�@N���!�Z(N��g�V�u��y���\_m|Y�n.�7�m3T� ����@�>՟�U�{��@;��g����K%�����Uũ�M_��b4��2Эp��v�Kv��n~�:��l ��&�	��mf���P����1�o�2WE�⍼���RR`�i+\(\�/{��#�*�|ȉ<�vk���'�N�W�S�7z����~3���qj��Û=���"`�NGA�TQ�u�[!B����nk�2�e	t�V҇�l����~�Q���MFp���)�>�4M��g���|t�@_xN�ѽ=�x���f�*�}P�s�T�a���pTb��#4�Cj������5�q�e١�@ ��C���V��բ� 7�:<HU2�g�Vl��V���e���j����&c�Ql2�4�n�Э��R����T�9�us��$5ށ^!��3�!:�O�
��nbJ��OY6���F��2�MMN,O7�᫔�W��H\�}1�:����_���7�w����eGR�f.���/�(���Կ�&��g�k��&�z����Iی���s�������1j��^�"���g<����c�	r�/)
%Q��-ۼ�,�Bk��9�z�}T����7��e%o��f��Cb�J����vZI�Q�%��|FQ�$�)C�n.72��v�I<�����s�#pM<V:�R �,�m.�b�[+qc��Ǌ/���\x�Q'�+?ƍ��m�/݂8������8�,�U	�ۭ-e�o2���l%�����r !N�ݢ��/��zi�6��9Y�J�V������Q6����i�X�B�����ݶD>�<��#x�I�.z#���{n�!��0]#���[#����J�q�S-]�NY��+ƍ�=�����is�8��U�BZE�3쮉_������8!�6��j�z'~iO��N�^����a�Ɠ�&�BNAm��B���O��m����8�P�8V!�`´lS�a|w?�%i+�#\�����[��2�Πj�v�E��&�i�nd��i�Y���c`��lh�!O1Q<n$Bޘ_������-�"�qk)}3�Ή�V�7���H�
ĕH�	�t�%�Y ��$i� c����Ėx�܏񨨥,Iϋ# �V�l%����Υ_�p�p߉�=e9Q_�E���uhf�>o�d��;��l�~�� �b��ߏ���ƌ�ST�}H+�˾�'�S�i�s����渉_�<������%(l��z�K���ɋ�C�Hw� ��y��+� ��|樂?}d�)c�܄/[���5��;�X��@1�Vڞ�P�"���N2+��7A�v��4Fx��J��P�t%[�^4�M���j*�N〉L�=*ٍǨ]�zD�8�>���*�J�D�?�~b�9����R����劔[~ᾐ�O�E�R&�M���E����\�������R��(��p��������c�DSJx��y�G�`��Jˆ ��G�r�ܯr|*�P��S�:e�3�^��1�m��g��6%�~1(��U��z����E>�eS9�r6�n��)lX�W���U�(����jb�6䵥�qN>���~�U��֞�zQ���5�o����!�fz�H\�Oz�OT�S"���z�����W�o���l���2H)?��jg �5�`K����Xց
��z���QZ/z���J�e1	v7.-DAM}F	�o��L��&��q��gc�04�� �C��0*���,ltl�K�X[�Y~_��O����_��	M7.�KL��F�ҽ����E��C�������,���.!ߛ�7|�	@n�l�'͍�e��`h�+�ŀ��)�C=/�th�}+����3��(� �2Øg�mO�L�t���?X����h ��̷�ע�?��n�
�خdH�j?��v��Ĉ��
r��آ��2}���`���)��Z࣐���B�P+"̝V�N8����zu������Jѯn>�̒����W
�kf�����k���\�g�yK+R��i&!�l��Ξ�"�$o7�����G��_���O�A���-��6�R֧4u�wa�)o��,A�3Ͼ�M��9�5/c+��x�7t|�8���ԯXr��0��=X# �����|�C~r� F�� �!�ۏ:���O��E�����GT�g���m� ���D>�gR-@S0��Z�d�褶t)��j��}3A(&J�'�O�'�����՞D�Ñйo�i����N++��g(c�ˢMh���5����
[>�F��Tu-��)E�bCZ�=���ɛ�O�����, Y.�`�1W�:w��^ٽnO�%D��W�PF{<�+U,��O���cd���OX��=����Bk-"TpI��� ����Y5jN
Z��&>��燯�hWC/�ۇ��@-z��w��D�6�kOЫ����_��M`9��8h��iCX�� ��L
k�͏�>��z��,jɌ����{���g��l��f�{ h�Zӈ�^��|k��v�J�����@�ʠ�h/ .��u)��׎����L+�x�3��c=i������G����a�7P�ew`X[����5W��q� ����]��Z�9�R��r^����c�xz����~|i�: ��"6c��$��z�_�?nQ�J���T�`���9"S.M��nQ�^R8E,}B��iR��ڨ<g=�����
>ɲ���p��eO�ͩb�v�U)��h����[�VB�2�e����K*LJ�/�]�J+Ux���vn���H��4��������m8uС ��\���؋B�Xy4���r��:�U�5RE��>����β�Z�uш�jUz�J�w A�@jDm�n��6[}}h����*�2���~�x����B">cN̏l0�Vu�Y��C'�y�IK�8��W�(�{|$���N���mܛ{B0:Z�?:oǞA��eFr�2���ڭJ� ���ado ڂ��,�l�l9y6�s>I���O<Κ��dP\����I����E\U�gn�YC ��d�� �DS���3;{�{�s�Њ��$�׍��tAf��p��*�fzG<���6������κ]�[�~%F����/�£��>�ɀ��@�'���k��G�,~�HlH���[`��VNC�֋c��$�>*�l�C#�*��?$����tY��_�G&���Q���ޢ;���^=|�}��	�U�j�W^b���l�y~f|�������"�ZT"?���O1_���8iE&@���/��tu��s��i��eL,���̕�U�)�e�k+1�3Ï{y�:<�#��3��S1���ߍ�Y��]���V���O�Ѳ�T
[O1��.��^~~��"�;}�F�r�g��D��kW�֌�Q�~��I;w��xf"��3u_��d�҆�&�մKn{w�+ޡ�B͕�K�0���*����=�;Qg��H,�@�$Ѽ��o��⪼G˹ZjQt��b1��1�d��t�!�d�)3�=��̗kB-���t(}2�A�G�GƎ&�_\T9�P|Ҩ�<-���WhӀ�.�B��oepR��t����:��ũF 0���.e��~(a�7�e��J�e*w?w�yjR�-���X�0��P6#��:�K�-6�6>��+b���K������(2��l"Z^�,����/߲G3��<��ٸ���a�Y�|� ���"M����ۢ��xqd�E���J��`3h�!#1{��ۚ�:���z����<�^���R[m4�{����y�[�E��&dN�s���>a���S���AD5Y�����K��dah~ K��k�4����F����{#m�����i5��ad���3L
����V!��g�+�P�`��#{�gPaI)Q�.o���M�d=U�q�
�Q�,\���>�"�`W�h�K.L;��5��'�� ]��b �S|gQ���XC_����iMa�Q	�4ծ���P���Ȉ�g�GSkI�	$%��c��Bi[z����Ƣ��_� �Bo����m�ꅷ�Ǩ� 3PPН���F}����]߀U�qV�n=8k-��c�;L�7	K�{����_
��l�>���փ�B=m��]A�т' &ˠ�':�(��y�d8�e3���.��0�Z�|��	^rN���3��~5ǔwzru7W)�����g^�d��5	�B����h��eIj?G���b�/�����͇�[R���h��'p���u��.(L��P�Y�rz��~��KKX��f:gLKÎ����U��Sm"���/Y�-���=��#8����u+��H��Rݘ��P�����?��!r�79u�6e�)*�����k[�;��X=J�J��S�>�>7�����1��f���[��s+x�G�A�9�b�
t�>[��@�`8���/l�]'t۱rŕWKK�v�ڙRE����
|rn�º����5�n/$����|�=@((a���=mO��	�>��cYa1I��O�TO����T��Ύⓓ49`���*e��	̨���x�rZ�8��Ov��p�����O�H뷔_��yn���-m$�J=�`��7�V���F��g���pm!����փ�A�lй��\�IPn9�i!�:�߫MR�I53��f�	�uu�$����/��O�0� �Y1U���6�
ꔯ�4�5D����(��w��}�t/=| [�[�t���I���_����h�s1x���N�
��]x��Y<����½�1M����Q��(�S��Ɏe�2ٸ�D>���Wtp�*9�K��P��Qt�\BC�'�й^Ʊ:ʓ�M��3�9S���pr���ܵ/0�뛦�z�;w-��������__�(��1cR�%D��r�-k�荼�;s��ݏ'~"wH)��I��r�]n�a�ȣ+��C�����n���\*;�G��q�͏��d����1�~�����s�,��m>�P �ٶ��c�j*}�G�!	�P�?����M�aS��K|�
HeM�{3l�<���:�7'�m�a��ϛE��i;��iC!QK:��t�׳S>�8H�{��9d_�.���N)I*Z��l�YA)�6��QS��6f�;l1�~F��3A���|9�n7���s��&9-�����Z��л,[�4Nɯ@��<��#�����'+���X���]�����f�?U�3����[s^�	��ֈuW�z���4�#Ҏ������E�/�u�W��;��:�������a���2�)�!2�9�Re��g��ô�d��vSߝ0w�zbg�B��_�(y��H�$	��A�#wD*��f����80r��!����+
�~�D�U��Nגh�A�����)Uݏ�S��x���@I�'�,��f�W_�TZ�P.J��2Ɲb�Z:��/�^G�� nyH�!��"�VM>`��ѧd��^_)���ny�;���~�
�O�o�!��N�ۗ�C%��Q��U	��72ja����1]�O%CLAY�WI�}z���鯦���	$J����i����lO�^#�^q]�a��_��T�m�2�ک=���a��G`�hn Z�MG��u�ϙr��ny�h4�z��bMJX��1�?Ň��*�Mߤ87#��}���ۖ��MD�Z�x��D�����K��<�,���5If��X�O+�+��G���q ���{�B�e�*���[SbY�ź0dϒ� ����Ɠ�ɿ��K����:��B�"�r,��6���X	s�IY-�d~(ɦ��jʇ�Cй[T{�EW�2��o ��d~��$�ơ��;��j~�B0����S4���J�J����S��h�'���c{���e�ˢ"���c�p�(��Ô�ǿ��������]�� �yp��K�c�aGc��GU+4I>����h��^�x�NzZ9�O�k4<��~�t����[�`،����u��D�,˹�s���l��	\ �1J�x���f>_��+��hDdí}2�Um&���}��i�bxW���D[�w`��W�7����p�D����~�
Φ���	ʬ_BhH�4<a����9�+�d�0�*6ds�a؀b��g=|��XhS_) <r�T�Ɂ�@��ǳ�[K��
�2�#qܗ|��@����^�����7�a��sȫ�
�f�c�R��e�
LAe�Ԅo��v�����=��P1��j�nI�t9LsY�I3r��S�&�r����@�=�O��r�3�i�l�RBK��ևZ/D��0$%4�<���v�ۚe%3�D�ӛ �:R>1��+���;v�x.?�a�'�(����s�����%�R�h�XJI��ا�3�$���z���;J̫Hpל�z� x����>�V��Z�_�om��(r���ve��]��2(@��گ�L%����l���EM���Ys]1���O��B�_��(.�D���ʬ'f��Y17u�$�+7dL�~yyf�N���c<l�i���Rd��:�k�a�"}�ﭞ�Xߥ�Q
�$pKx�������	���X{�VI�uMP����Þ<2r,��)��Ѧ�l���ʦ�n�.؅�}�I���B1����2�\����c��`K\+>�s3l1_�w����6���F��h1�h��9�_=zgO��q�Q1.	�#l�~P*ir�\G/f~�}���3DĂ46$��9�

޻��϶�ر;��a[#�0�$�Q7 *ˉ||�M1,h`�	��N۟��0��BO���I�uI����$�V*\��f�'h�H����]S%��� �C3o���o�+�p�(�}�~*��S�񢛼��K$�
�o����%[��,s>[T}��S��ޏ�Ǘ��3���d�ڿ��
0pV�j�cU_�W�d`Q ���d8n�07�lȫ�P+�P�V5����*������J��6h;0}��E���+���$�R"ߨ�@F8R�${�K͟��4rm�5Em�@`XL���d%�����a��H��km=�B�d�Mt��a� �Tf/^�>8v4ƅ�U��{Ͽ��?s����B�����K#�L�'�hT�^~j,�nu�������ǁ��C���j�U�PI��JGx�qݑl�;��U�4{A�Ҁ}tl�HiɌ�W�=Y�M��˧)m�@�~��r����0�r]�w�^S����WU�p�,L��YZ�q4Ec>t���(��@�C���o�z��N�l�oz�V���L8�3�APЍ�����I4�j��}k���̤m.��jDȓ�l����H�v�^XjS�X[,���S�~��6@����:Ɓ[��y�h��r�;<�X/:3�ܙYZו���\>s^�C���<�J����"^^��H���q�M<�����߾��7Z^^C9+g�I�6_	�(����u���}H��ԣDiz�f��o��Hr#B�IO�ya�2��ַ7$��J��ana9$�V��k��wŋ�m	���[���'�8�H��G���\��0�TJ��I���r�}/ l�>�m~���'�\L:��1�61�]�ai����W���i� D��k|t��x�O��uMJ0$ߌU���BW"�z̸�c1�M!ͼ��K��胁����^��L�&��Uc���&�;Tn�;\�����i�fj��� �j�8�\����#XV��d{a�m�J��q���sk�ʹ����n��	A-SN���-����v�?��%_�us�:2[*��(pQZ���1����;�[q���,����┄�#�� ��@��9Yφ9�W�g��˟*Y�|��QT]^^��H[�1A7�&I+�qx�����	SX��D�e�+=A&�;�Fu�}�]J���V�Y�g��t����Vs�=��@��/�֔W�x;f��gt`�����
�3=����5v]Kv�m��H���O*"}���L�l$�;��p@�����h�괺�B�Vvn!-�4�4�4A�ոJ�����P(�kwѱ�Ak��\����h��8{t�2sK�� ���	Vy?�~?�:d�l�CQ��]\��E�B��L�����+F"ܮW� #����yA�j}�1p����,c�7�-vA
��8�t����ܪǾd}�O�Z�������'�����zN00.�'�V������FXrǐG;r��1y/O�B�|���������6���*�.�\�w�[�Wr��S�`É���5>X�< ��SԞ��,~_���5,�|�C^����7Q���T��4�J 5���m���q����R�����'�[���ϸT�U�w� ������+���{a�^U���y;O����~��od_��2��d�Rg~pX�O�e����+v����=<�4�_�Z��Վ͝�=���$"�Z��Ir۟���>����$"�,�3�VǷ�c����++uK�-��PgW%e����\ꮮV�U�=����J7ϯ�Q��_׮��Z�T�ё���D� ������ji75�0�U�Z�v}��h>(UW1yG��9�6�꣰���.Ȟ�G�r����[�sn��#��	�Y�i�@ޒlx��}G�
�#��m��$w>���?� �ɗ��0\Qj��S��ʔ�#_�Q\ �x��e#̆6O�Z�l�i��a+�xKV�K��7!�C��Х�X�~v5|Kb�(�����0�/?/��W��׏�%ߴ0��8�hV�v����	K�q$R��T��x�)���� ��i8�q�Z��G.~�:3NmV�
nB\�����c���$�!�D�����	�rEi t(<t6��3���.�~�"��nP�.���poD3��lp�^��3�;�;�"�z9�3Y
A�i7(n����}=��>�>�b����t�P7�D���f�]Y;ׅ�
�]�l��=���t@��/B��z��K5��U�va�?�ov؃o��ZbB'0�$���4��L��V>b�`Z1�ވ��S0�j�J��`{�.wvqKӚ��M@����@?fc��6�@��c^���ewÌn
3\3p-�_}ui��!^���Z8���l`O��"<���'m��?g�l��n��6�Pg�"��|�6��ʡb���Ig�I�O**clnOV4j�vD�Cn���]o"����ۜ����(k�O8������oz���#d�h�|$i�~g2���)������Hb�h�h.i\*g�[���o�B�_R�iMKJ><��̏R�1�ŷgB0!�F;>Gڶ!-j�b[�	^�Dz�F�<7?�-B{��T�c��
�*l6�wYz�	��K��l�4�c;Cj�v�}�'�����7����5͆�.���W?�����a&���ں5��23@!z{u����_��^?J8�4f�wt@��2�sP�ʩp��%D�Z�_I\u�re����<if9�h��^��"��x��� pX�����>�M�g����,|����]
'�h>�pr���n	�%υ( -q� ��e&�K���O�����a9} �q4���:����YVE�;��@e/2v��3�U+�C���c�Kv�Z��r��vR��װ�EU�x�xLkSQ�:-4<0Q�W� �M$0͐�H�+�x �%Ák!/Gv2��@6A}vE���|��(�U�K���>��;"����A������|_��e�id�^
?��*i#�V��\�7�?�n�0p�O��	�_��Q�(�Z�ޝ��9�/2[C���bB2�����RN2�M��U#���)�e]M gZmn+�(T�L{��z@+�.��s��F������D���C�q��5�KG�R�UX8��OB�ѭ@3!�ИB���}��K5~������!���V��mG�`#�� �Df�l)�L`V�Ի���2q�����[c���7X�/�v�`w8����ƣ���Dy�*0���oH�
���^����)>�&[D�cf3���� ��Fx|{i���C����N*49ɫ�eN����;�ȳ²�^?8�ڣ"��:zx���.�!-�`���z�n� �z�#8+rN�����Uǎ�qI��g���0���q�@����"0��P��"���
�^Ɍ�����Ý�E�Щ=ߣAPp�g_9I�^R���]kg����$@���tJ��-����_��I������e
�ǵ>*D=l��k��'�s��S(Ġl�A=����QC�6w/����x��	��p�9�/��7���=aP�?��s~{�/�Mޜ�,K�Q��h�nq~2���!�מ/�\��)�����.G%���z@(��1ʖ��7�2-�t`@��6�B�n�Jt9��:�7Ly�5W`��T�d-����q�͡�����Y�^Ӻ~e�c�ʣt��L�p��Eо_wT�f�o�r\�27Bt£8�n�T0Rs;h9ְ�U�3R���Y8]���� <"|v8��q���+��B��?�(�Q���}s�r
�\o!�ץ������[W�d�u�Q4�Y�FQ�&D)R�w:���⎭��ʾ~z%\� ��ŗ(�-�]v"c����S��wu�e�:��چ���� �Z1לJhj@�]����9�V/*��J.�����7l#�i�_�E$9��3M屯�q� �����e�NMxƆ�@���E�M����@'H	[����a���ʀ2�è�UX�~�=�V� U���/�8n�_����~V���Ót�/�a��L7�!���������)�r 8�����9�_b�󿬘�_\.� 
��?� �7
3���b����ཚ"!��C�E��pw|����'�Rj�U-_����N�K�.����y%�U�M�KcZ��Y�^ ^Q����$VЫ���v�)�O�r_"ܠ�&�$���u��0�])�Wމ�´������eT|z�����r�x�n=QC�G�;�����ʰix�-
I��ܫHa�bA������P�Pܼ��S�������LD�a,�" ��'�(��ޠa*y�����1�(M~�f��8�ݎ��!i��6մ\u��QE�-7߅��߇��սv���eb��8��|Z�>0�n`x�Ƹ�*W��Ț5�� �ͳpl�9D��2����鵯
�Bt=�����kU�ȿp��
/��O�������͖�~O���2֏��ըYW6�O�(ԹD���3��兯���n*a�j��Z�.��# ]��
���mC�S�&����Y#ƅ�f ��Q�Ds
�v����>C�.���:zK몌=�ɮD�xn�3�o+�l<�H?q�噄2 >��i��D�`3u-e��R6<�d�i�@pI�\����Y�o����>ǩ��_�5�H:jlk_���f�N:hA��Ӡ:Z��;(�3+b� A���"��<j�h��m����{ ��P�sx�H=���Ԣ'`�7�.{�h˹�ȅ�"+s���)�E`%��͸�w\0չ��n�:o�dd��5�XA\c��7�K����t���/���e���8�O�ꢂ����8�)�5�����]i����b���G{eW�5�0#gP���GM���5���]���`���2b�c;��
`��$���ҽ �Ս�)����<g�ߗ�V��ѓ����D�
����g[R�c<zZ�I(i�E����\b\�1r?Yc�����1�3��mߔo5
���zMd6HT��ޖKF�K�(!îAz�^%�M]��#��]��6�M�'.���3"���;R$_A	6�Z8��Ƣ�2H�gq�IQ�c�V�����+k�������7X =T�)��j�E �U�f��yWD�|�1|4<�_>�; (/~��<mcT �=$��D��w�@E�I�}�����?Lp[{c����5�-�N�Z3;x�z{B��,�����|�{gT�:��pȋ�Y�t�K���T"&�%YJ)q	���ύ�lM�1�G.Y�M6�%`L�a����J9��1�M�"�3҈�����V� "U�ݬ�<Z���_�q��{5�~��x��ߏ�UO����*��Ã0�Y���@D] �7N��B�rI�N��Ib��y�7�)v?��q9���ڃ��,Kfs��^�ೀc��<�6��$b	��kR���ȿ�NK�����������9�rz_�����:M��a-�\m��f*�>�qh���8��t>I��Ŏ�گ� 9��m���
�� �x
d����R��K������p[�yKy�;���l����Ď!X/��+kK�~~�_i�Xk���&�o_�E���n��fNf��#Kdy���I*��#�yg`�萣�sޠ5�F�R�N��jg�W�nu�Gc	>%��8L����`��K� �Wӹye,Cj��&ּ�u�*�^=WcY3_h̹��Dn�8� 'q�z �����m1�<��ڼK�ً%m��/���U�/L��U�-�kXS��{ J(#9��i*��ܻ`��=.�a��c�!~�p~���_��ܗ�I��5��do��(�8�ɚoC֏b$��y�$�<:����񜏝p_��H��o�K����(޳']Seh�jf{B�Nr�9����QPR1��R�ډ�!�-���*�xo�Mc����p�V�����oS�ƨXZ�Q�볂ȉ6�yRj���B�<�ci�8�g-}����a���4��ڄ�J|]ز�(h�s��ɔMAjO���g?�l!X�u�d݀��T�|���H�af#�y�%�u	�D$ yC�
�*�.t �RU$���pH�l�����|R�x�#��Ly(��e��������r�`*@r���wyl�ݔ�L^�L�Г��7��(-��Q�'U6�7D�B��MN���-o�/4�j�H�_?�(��e�o���U�	����s0��D&>�hh� ������J�&��0�o�3��<���.�3��[��6�mȨNMs�jjZ��z-#��똙������_AO�jot�ϱ�`n������ͻ�r#�}�5X� P������$�$����N�Lo��{�rmr��������>r�Ł�[�ѪFQ���i�`jL������:8O���e�k��I�P����E���C�q�*z�,�����`$}>i��3bA�?F���߅yy:ݞ�Ł� H3��Td~��yL�;괫�
 ���ǈ<�n�}�j��兒�Q���vBp�ۙ"�y�S�u��sR��o�|Y\�P-�����^�m���1��9'_.�C:Y�A��,ik��(���f���]�"�p��*+\�7j��+��/\�W_������|W�[�'c��u�ZpG��!ę�-R&M$q.��� ׫W��۔�+#�5�1�i�P��ǥ�X��nQDW�(K]�F:�E�YS���[���=M49Uә�C<{��l`0�	~�N;ƥH14:��"R��*0y�V#�*hܑ�J�S�A;��>3 �W���ET��xB���f�̿|&Ûk�ɟ��0F��Ƿ�J�P�hn��T�Ŝ@���K[���Ӷ �r�=<4T�S���u=�.�d��=�UA�}I�P�{)v2�M����	���r�x���	Y�x���o���jV����W̺���(�7�i�F�@�/���]����3����W���H�'��-��.�*�r���� X�l��������s�<�Ɠ@��v �;T�@J��ļ���o��$I���e_x>B���@�E?l����Ͳ��~,���M��r��.���No�&;a�n���*3�2,�!��m���Nė����Z~/6ޫ<.�M��"��O3���+�S�sl�/yir���<��Ou�L�,����Yl��q=����H�@��~�X&(� �E�J����t���!�;�C&fF�zsc=#�JT�S	����Q"�*Ф.6�>���_�ܹ%t�&xq�&�0Gܪ���Z)�`��$~��l�&W	�a�(h��5 ��N�@�I(I����B뱂�ׯQ��xN���pΦ�煟J7�Ԟ���� ��065�a�˿_��ඇ#*s��g ��IL��G)��{����$����Ќ�O�k��";a�@�n�~�sW꼙�u����#��[���K���yMPd7�OW)l��d��s=ԛ�ֻ�O�����X 2M2��A����w��%σm'4u�o��_}%0��l2@�ߝ�p��:��R��M\���Ι0��U�K���OXYǍrT�4�T�x����9~�6��hQ@ju�s���D0��Dp#J��3�*��q-��8>���2��.�k�{����Ÿ���}`�e��d~�bҮ�Ӑ�10P��/'j��-1�eF.���%����Gg�����1+�z��
|���d��nl�ν�[XK��E&��V�������a5�Q9:��m�Qc��U*O./+�}��"�G���[�D�qFE�y)^�m��^�:뮨��f&0�i�^�X�g��P�H���^�6�	�>Q�ۏ��=�zF�!x��%[O�7�rQ�L��K����ޥ@��kɗ誗�{z��'�Ϝ�d@�!L�@�E,����Q�+�S��'{f.��Fr�)���8nf]�c�ܡ}�zVb�4����ؖLi���������8��\��N�Z��	H�-�9����*(QX�%c.q� ��l�W�HF�4<(�6OXmp�����/jW�8�Fu�H��QYS�rʻ������e���pC`Rl���[ ��	v!�Щ��
JݵF5�2-.7�Xs�bi�o��Ml����N�mh�;<?8���r��T�L��vn.Y er,�jA����p�Z��
����B�מ��D�0�/�&\%�%�&l�ܠy�D-vr�:�n�q%��%]Ы��7#���4��z!�RR7�حh0D>�zs�v����	�q���l�"~^����(I�F�!���nZ���[�����l���B��w��(u1����NE��>*Tc
���-��>`U%���׌2���B�cm���
�;�O �J��4��_g��Ӹ��z@�9JB<�v���(��i4; .%io�ב�%�b�#�"X�[�HKz�ۈ'��R�A�-�h������}:���mL�^�z��70뗨DCDp�@%Eaq�YJ��㒑�K�o��1�wؾc��3:6� ��"�a�(�b^�i� 7y�� X&^}p��w(¤�=�-8b��ĄI�uw�]�/ݠ]����{��]�(4+�-�s�\�,� ��e���H��V�[�%/����Xun1�2��I@;jW(h!�#���������q�LƼ&`�a5��~O��/g�Yj
����%�_�F�KK��a3�#�Mc��9�����'` ��'�|�f�H�$��	�_�\si���hV]����=���T/G�9��&�Tf�A3&�ܰP2^�&�SI������$��zu� �1\�H3-$-�u%�{��~����ٮ�\���L��+���9Z[4q�܈��C���/���KQj�g:@�+��ZӔ�c��y��sZ���2��蚟}��[�@g���	���+�v�����5{��`i&P�C�JQ��q��˝r��
����h�XN@���"ļɬ����V%f���7^<�j�bUF�\.�U�$�0Ԕ	�m4�f����m�T�~m�ą�*��GfC��u��������é���Xo��f#�! Ӹ���o�:�'�S%��_feN�
�Ď�)��?ov�E� �r}JwQH]wJ ͻ��틙=���|�R�8H�Vcf�)K]l�p��Z�d� y˦��Y�p�k�څ�f��L�b�3�
���u�K,�>B���?�*M؃��5�b@k)Φ��L�L�����7���IAA��iW��G����|�^��,J�����%��ŭ�v�W��4�H"
b$�2�W���FM^��0��|�DG�<FD~��Y1|܊-����+C]�&�"��0^�);VI��os��B�L�[q�������Z�סD�N����J�8g��vi��Dftq���R�	�y(�t���/�wM�~�(�$�S����Z-��������0U�H��1aolwcV���"&l&N�V*�<�`D�q �e�o[M?(���X������M~#����i���һ�H^���vEJ��+� �뷈�Ts#��g;�w���C�N���!�<��	��TdmV���!���5�!��[����w��4�iFhq�I�6���0�[|�D��&3n}��CD�Q�a��,�R�3���_�f��8���"�����Q� ���'��ΘYN��B\!rج{�6H���u�T9�K��/�Փ�Hڄ� 'S8�����/�� �+�Q�.���~��t����d��6�Ϳ	���N(k#�u�������^唕=������m�p�ُ�j{�~��#g9'�&4qn�#�M��.��z�;'����8�W=����53;�1�wP/�}@V�T���0e{����͍�
X�z�:�!�8B�mt��y]uE�7{��ї�;��u_!l�P$�7�d��H�	l���;�ϋ��k�&��o�X�WbNÞ�T+e�q/>�P�q|�S1p]����/p��͂e�<0'���� ����	�	|�|��^��,앵V��_�3�ʆ�����D���(��ى�duQPA�
@��Qs-�jK{a�g�